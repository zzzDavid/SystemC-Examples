`timescale 1ps / 1ps
module dut_Add3Mul2u29u8Mul2u8u8Mul2u8u8_4(
          in6,
          in5,
          in4,
          in3,
          in2,
          in1,
          out1,
          clk
);
   input [7:0] in6;
   input [7:0] in5;
   input [7:0] in4;
   input [7:0] in3;
   input [7:0] in2;
   input [28:0] in1;
   output [31:0] out1;
   input clk;
wire csa_tree_add_48_2_groupi_n_0, csa_tree_add_48_2_groupi_n_1,
     csa_tree_add_48_2_groupi_n_2, csa_tree_add_48_2_groupi_n_3,
     csa_tree_add_48_2_groupi_n_4, csa_tree_add_48_2_groupi_n_5,
     csa_tree_add_48_2_groupi_n_6, csa_tree_add_48_2_groupi_n_7,
     csa_tree_add_48_2_groupi_n_8, csa_tree_add_48_2_groupi_n_9,
     csa_tree_add_48_2_groupi_n_10, csa_tree_add_48_2_groupi_n_11,
     csa_tree_add_48_2_groupi_n_12, csa_tree_add_48_2_groupi_n_13,
     csa_tree_add_48_2_groupi_n_14, csa_tree_add_48_2_groupi_n_15,
     csa_tree_add_48_2_groupi_n_16, csa_tree_add_48_2_groupi_n_17,
     csa_tree_add_48_2_groupi_n_18, csa_tree_add_48_2_groupi_n_19,
     csa_tree_add_48_2_groupi_n_20, csa_tree_add_48_2_groupi_n_21,
     csa_tree_add_48_2_groupi_n_22, csa_tree_add_48_2_groupi_n_23,
     csa_tree_add_48_2_groupi_n_24, csa_tree_add_48_2_groupi_n_25,
     csa_tree_add_48_2_groupi_n_26, csa_tree_add_48_2_groupi_n_27,
     csa_tree_add_48_2_groupi_n_28, csa_tree_add_48_2_groupi_n_29,
     csa_tree_add_48_2_groupi_n_30, csa_tree_add_48_2_groupi_n_31,
     csa_tree_add_48_2_groupi_n_35, csa_tree_add_48_2_groupi_n_37,
     csa_tree_add_48_2_groupi_n_38, csa_tree_add_48_2_groupi_n_39,
     csa_tree_add_48_2_groupi_n_40, csa_tree_add_48_2_groupi_n_41,
     csa_tree_add_48_2_groupi_n_43, csa_tree_add_48_2_groupi_n_44,
     csa_tree_add_48_2_groupi_n_45, csa_tree_add_48_2_groupi_n_46,
     csa_tree_add_48_2_groupi_n_49, csa_tree_add_48_2_groupi_n_50,
     csa_tree_add_48_2_groupi_n_51, csa_tree_add_48_2_groupi_n_52,
     csa_tree_add_48_2_groupi_n_53, csa_tree_add_48_2_groupi_n_55,
     csa_tree_add_48_2_groupi_n_60, csa_tree_add_48_2_groupi_n_61,
     csa_tree_add_48_2_groupi_n_62, csa_tree_add_48_2_groupi_n_64,
     csa_tree_add_48_2_groupi_n_65, csa_tree_add_48_2_groupi_n_70,
     csa_tree_add_48_2_groupi_n_71, csa_tree_add_48_2_groupi_n_72,
     csa_tree_add_48_2_groupi_n_73, csa_tree_add_48_2_groupi_n_74,
     csa_tree_add_48_2_groupi_n_75, csa_tree_add_48_2_groupi_n_76,
     csa_tree_add_48_2_groupi_n_77, csa_tree_add_48_2_groupi_n_78,
     csa_tree_add_48_2_groupi_n_79, csa_tree_add_48_2_groupi_n_81,
     csa_tree_add_48_2_groupi_n_82, csa_tree_add_48_2_groupi_n_83,
     csa_tree_add_48_2_groupi_n_84, csa_tree_add_48_2_groupi_n_85,
     csa_tree_add_48_2_groupi_n_86, csa_tree_add_48_2_groupi_n_87,
     csa_tree_add_48_2_groupi_n_88, csa_tree_add_48_2_groupi_n_89,
     csa_tree_add_48_2_groupi_n_90, csa_tree_add_48_2_groupi_n_91,
     csa_tree_add_48_2_groupi_n_92, csa_tree_add_48_2_groupi_n_93,
     csa_tree_add_48_2_groupi_n_95, csa_tree_add_48_2_groupi_n_96,
     csa_tree_add_48_2_groupi_n_97, csa_tree_add_48_2_groupi_n_99,
     csa_tree_add_48_2_groupi_n_100, csa_tree_add_48_2_groupi_n_101,
     csa_tree_add_48_2_groupi_n_103, csa_tree_add_48_2_groupi_n_104,
     csa_tree_add_48_2_groupi_n_106, csa_tree_add_48_2_groupi_n_107,
     csa_tree_add_48_2_groupi_n_109, csa_tree_add_48_2_groupi_n_110,
     csa_tree_add_48_2_groupi_n_111, csa_tree_add_48_2_groupi_n_112,
     csa_tree_add_48_2_groupi_n_113, csa_tree_add_48_2_groupi_n_114,
     csa_tree_add_48_2_groupi_n_115, csa_tree_add_48_2_groupi_n_117,
     csa_tree_add_48_2_groupi_n_118, csa_tree_add_48_2_groupi_n_119,
     csa_tree_add_48_2_groupi_n_120, csa_tree_add_48_2_groupi_n_121,
     csa_tree_add_48_2_groupi_n_122, csa_tree_add_48_2_groupi_n_123,
     csa_tree_add_48_2_groupi_n_124, csa_tree_add_48_2_groupi_n_125,
     csa_tree_add_48_2_groupi_n_126, csa_tree_add_48_2_groupi_n_128,
     csa_tree_add_48_2_groupi_n_129, csa_tree_add_48_2_groupi_n_130,
     csa_tree_add_48_2_groupi_n_131, csa_tree_add_48_2_groupi_n_132,
     csa_tree_add_48_2_groupi_n_133, csa_tree_add_48_2_groupi_n_134,
     csa_tree_add_48_2_groupi_n_135, csa_tree_add_48_2_groupi_n_136,
     csa_tree_add_48_2_groupi_n_137, csa_tree_add_48_2_groupi_n_138,
     csa_tree_add_48_2_groupi_n_139, csa_tree_add_48_2_groupi_n_140,
     csa_tree_add_48_2_groupi_n_141, csa_tree_add_48_2_groupi_n_142,
     csa_tree_add_48_2_groupi_n_143, csa_tree_add_48_2_groupi_n_144,
     csa_tree_add_48_2_groupi_n_145, csa_tree_add_48_2_groupi_n_146,
     csa_tree_add_48_2_groupi_n_147, csa_tree_add_48_2_groupi_n_148,
     csa_tree_add_48_2_groupi_n_149, csa_tree_add_48_2_groupi_n_150,
     csa_tree_add_48_2_groupi_n_151, csa_tree_add_48_2_groupi_n_152,
     csa_tree_add_48_2_groupi_n_153, csa_tree_add_48_2_groupi_n_154,
     csa_tree_add_48_2_groupi_n_155, csa_tree_add_48_2_groupi_n_156,
     csa_tree_add_48_2_groupi_n_157, csa_tree_add_48_2_groupi_n_158,
     csa_tree_add_48_2_groupi_n_159, csa_tree_add_48_2_groupi_n_160,
     csa_tree_add_48_2_groupi_n_161, csa_tree_add_48_2_groupi_n_162,
     csa_tree_add_48_2_groupi_n_163, csa_tree_add_48_2_groupi_n_164,
     csa_tree_add_48_2_groupi_n_165, csa_tree_add_48_2_groupi_n_166,
     csa_tree_add_48_2_groupi_n_167, csa_tree_add_48_2_groupi_n_168,
     csa_tree_add_48_2_groupi_n_169, csa_tree_add_48_2_groupi_n_170,
     csa_tree_add_48_2_groupi_n_171, csa_tree_add_48_2_groupi_n_172,
     csa_tree_add_48_2_groupi_n_173, csa_tree_add_48_2_groupi_n_174,
     csa_tree_add_48_2_groupi_n_175, csa_tree_add_48_2_groupi_n_176,
     csa_tree_add_48_2_groupi_n_177, csa_tree_add_48_2_groupi_n_178,
     csa_tree_add_48_2_groupi_n_179, csa_tree_add_48_2_groupi_n_180,
     csa_tree_add_48_2_groupi_n_181, csa_tree_add_48_2_groupi_n_182,
     csa_tree_add_48_2_groupi_n_183, csa_tree_add_48_2_groupi_n_184,
     csa_tree_add_48_2_groupi_n_185, csa_tree_add_48_2_groupi_n_186,
     csa_tree_add_48_2_groupi_n_187, csa_tree_add_48_2_groupi_n_188,
     csa_tree_add_48_2_groupi_n_189, csa_tree_add_48_2_groupi_n_190,
     csa_tree_add_48_2_groupi_n_191, csa_tree_add_48_2_groupi_n_192,
     csa_tree_add_48_2_groupi_n_193, csa_tree_add_48_2_groupi_n_194,
     csa_tree_add_48_2_groupi_n_195, csa_tree_add_48_2_groupi_n_196,
     csa_tree_add_48_2_groupi_n_197, csa_tree_add_48_2_groupi_n_198,
     csa_tree_add_48_2_groupi_n_199, csa_tree_add_48_2_groupi_n_200,
     csa_tree_add_48_2_groupi_n_201, csa_tree_add_48_2_groupi_n_202,
     csa_tree_add_48_2_groupi_n_203, csa_tree_add_48_2_groupi_n_204,
     csa_tree_add_48_2_groupi_n_205, csa_tree_add_48_2_groupi_n_206,
     csa_tree_add_48_2_groupi_n_207, csa_tree_add_48_2_groupi_n_208,
     csa_tree_add_48_2_groupi_n_209, csa_tree_add_48_2_groupi_n_210,
     csa_tree_add_48_2_groupi_n_211, csa_tree_add_48_2_groupi_n_216,
     csa_tree_add_48_2_groupi_n_219, csa_tree_add_48_2_groupi_n_220,
     csa_tree_add_48_2_groupi_n_221, csa_tree_add_48_2_groupi_n_222,
     csa_tree_add_48_2_groupi_n_223, csa_tree_add_48_2_groupi_n_224,
     csa_tree_add_48_2_groupi_n_225, csa_tree_add_48_2_groupi_n_226,
     csa_tree_add_48_2_groupi_n_227, csa_tree_add_48_2_groupi_n_228,
     csa_tree_add_48_2_groupi_n_229, csa_tree_add_48_2_groupi_n_230,
     csa_tree_add_48_2_groupi_n_231, csa_tree_add_48_2_groupi_n_232,
     csa_tree_add_48_2_groupi_n_233, csa_tree_add_48_2_groupi_n_234,
     csa_tree_add_48_2_groupi_n_235, csa_tree_add_48_2_groupi_n_236,
     csa_tree_add_48_2_groupi_n_237, csa_tree_add_48_2_groupi_n_238,
     csa_tree_add_48_2_groupi_n_239, csa_tree_add_48_2_groupi_n_240,
     csa_tree_add_48_2_groupi_n_241, csa_tree_add_48_2_groupi_n_242,
     csa_tree_add_48_2_groupi_n_243, csa_tree_add_48_2_groupi_n_244,
     csa_tree_add_48_2_groupi_n_245, csa_tree_add_48_2_groupi_n_246,
     csa_tree_add_48_2_groupi_n_247, csa_tree_add_48_2_groupi_n_248,
     csa_tree_add_48_2_groupi_n_249, csa_tree_add_48_2_groupi_n_250,
     csa_tree_add_48_2_groupi_n_251, csa_tree_add_48_2_groupi_n_252,
     csa_tree_add_48_2_groupi_n_253, csa_tree_add_48_2_groupi_n_254,
     csa_tree_add_48_2_groupi_n_255, csa_tree_add_48_2_groupi_n_256,
     csa_tree_add_48_2_groupi_n_257, csa_tree_add_48_2_groupi_n_258,
     csa_tree_add_48_2_groupi_n_259, csa_tree_add_48_2_groupi_n_260,
     csa_tree_add_48_2_groupi_n_261, csa_tree_add_48_2_groupi_n_262,
     csa_tree_add_48_2_groupi_n_263, csa_tree_add_48_2_groupi_n_264,
     csa_tree_add_48_2_groupi_n_265, csa_tree_add_48_2_groupi_n_266,
     csa_tree_add_48_2_groupi_n_267, csa_tree_add_48_2_groupi_n_268,
     csa_tree_add_48_2_groupi_n_269, csa_tree_add_48_2_groupi_n_270,
     csa_tree_add_48_2_groupi_n_271, csa_tree_add_48_2_groupi_n_272,
     csa_tree_add_48_2_groupi_n_273, csa_tree_add_48_2_groupi_n_274,
     csa_tree_add_48_2_groupi_n_275, csa_tree_add_48_2_groupi_n_276,
     csa_tree_add_48_2_groupi_n_277, csa_tree_add_48_2_groupi_n_278,
     csa_tree_add_48_2_groupi_n_279, csa_tree_add_48_2_groupi_n_280,
     csa_tree_add_48_2_groupi_n_281, csa_tree_add_48_2_groupi_n_282,
     csa_tree_add_48_2_groupi_n_283, csa_tree_add_48_2_groupi_n_284,
     csa_tree_add_48_2_groupi_n_285, csa_tree_add_48_2_groupi_n_286,
     csa_tree_add_48_2_groupi_n_287, csa_tree_add_48_2_groupi_n_288,
     csa_tree_add_48_2_groupi_n_289, csa_tree_add_48_2_groupi_n_290,
     csa_tree_add_48_2_groupi_n_291, csa_tree_add_48_2_groupi_n_292,
     csa_tree_add_48_2_groupi_n_293, csa_tree_add_48_2_groupi_n_294,
     csa_tree_add_48_2_groupi_n_295, csa_tree_add_48_2_groupi_n_296,
     csa_tree_add_48_2_groupi_n_297, csa_tree_add_48_2_groupi_n_298,
     csa_tree_add_48_2_groupi_n_299, csa_tree_add_48_2_groupi_n_300,
     csa_tree_add_48_2_groupi_n_301, csa_tree_add_48_2_groupi_n_302,
     csa_tree_add_48_2_groupi_n_303, csa_tree_add_48_2_groupi_n_304,
     csa_tree_add_48_2_groupi_n_305, csa_tree_add_48_2_groupi_n_306,
     csa_tree_add_48_2_groupi_n_307, csa_tree_add_48_2_groupi_n_308,
     csa_tree_add_48_2_groupi_n_309, csa_tree_add_48_2_groupi_n_310,
     csa_tree_add_48_2_groupi_n_311, csa_tree_add_48_2_groupi_n_312,
     csa_tree_add_48_2_groupi_n_313, csa_tree_add_48_2_groupi_n_314,
     csa_tree_add_48_2_groupi_n_315, csa_tree_add_48_2_groupi_n_316,
     csa_tree_add_48_2_groupi_n_317, csa_tree_add_48_2_groupi_n_318,
     csa_tree_add_48_2_groupi_n_319, csa_tree_add_48_2_groupi_n_320,
     csa_tree_add_48_2_groupi_n_321, csa_tree_add_48_2_groupi_n_322,
     csa_tree_add_48_2_groupi_n_323, csa_tree_add_48_2_groupi_n_324,
     csa_tree_add_48_2_groupi_n_325, csa_tree_add_48_2_groupi_n_326,
     csa_tree_add_48_2_groupi_n_327, csa_tree_add_48_2_groupi_n_328,
     csa_tree_add_48_2_groupi_n_329, csa_tree_add_48_2_groupi_n_330,
     csa_tree_add_48_2_groupi_n_331, csa_tree_add_48_2_groupi_n_332,
     csa_tree_add_48_2_groupi_n_333, csa_tree_add_48_2_groupi_n_334,
     csa_tree_add_48_2_groupi_n_335, csa_tree_add_48_2_groupi_n_336,
     csa_tree_add_48_2_groupi_n_337, csa_tree_add_48_2_groupi_n_338,
     csa_tree_add_48_2_groupi_n_339, csa_tree_add_48_2_groupi_n_340,
     csa_tree_add_48_2_groupi_n_341, csa_tree_add_48_2_groupi_n_342,
     csa_tree_add_48_2_groupi_n_343, csa_tree_add_48_2_groupi_n_344,
     csa_tree_add_48_2_groupi_n_345, csa_tree_add_48_2_groupi_n_346,
     csa_tree_add_48_2_groupi_n_347, csa_tree_add_48_2_groupi_n_348,
     csa_tree_add_48_2_groupi_n_349, csa_tree_add_48_2_groupi_n_350,
     csa_tree_add_48_2_groupi_n_351, csa_tree_add_48_2_groupi_n_352,
     csa_tree_add_48_2_groupi_n_353, csa_tree_add_48_2_groupi_n_354,
     csa_tree_add_48_2_groupi_n_355, csa_tree_add_48_2_groupi_n_356,
     csa_tree_add_48_2_groupi_n_357, csa_tree_add_48_2_groupi_n_358,
     csa_tree_add_48_2_groupi_n_359, csa_tree_add_48_2_groupi_n_360,
     csa_tree_add_48_2_groupi_n_361, csa_tree_add_48_2_groupi_n_362,
     csa_tree_add_48_2_groupi_n_363, csa_tree_add_48_2_groupi_n_364,
     csa_tree_add_48_2_groupi_n_365, csa_tree_add_48_2_groupi_n_366,
     csa_tree_add_48_2_groupi_n_367, csa_tree_add_48_2_groupi_n_368,
     csa_tree_add_48_2_groupi_n_369, csa_tree_add_48_2_groupi_n_370,
     csa_tree_add_48_2_groupi_n_371, csa_tree_add_48_2_groupi_n_372,
     csa_tree_add_48_2_groupi_n_373, csa_tree_add_48_2_groupi_n_374,
     csa_tree_add_48_2_groupi_n_375, csa_tree_add_48_2_groupi_n_376,
     csa_tree_add_48_2_groupi_n_377, csa_tree_add_48_2_groupi_n_378,
     csa_tree_add_48_2_groupi_n_379, csa_tree_add_48_2_groupi_n_380,
     csa_tree_add_48_2_groupi_n_381, csa_tree_add_48_2_groupi_n_382,
     csa_tree_add_48_2_groupi_n_383, csa_tree_add_48_2_groupi_n_384,
     csa_tree_add_48_2_groupi_n_385, csa_tree_add_48_2_groupi_n_386,
     csa_tree_add_48_2_groupi_n_387, csa_tree_add_48_2_groupi_n_388,
     csa_tree_add_48_2_groupi_n_389, csa_tree_add_48_2_groupi_n_390,
     csa_tree_add_48_2_groupi_n_391, csa_tree_add_48_2_groupi_n_392,
     csa_tree_add_48_2_groupi_n_393, csa_tree_add_48_2_groupi_n_394,
     csa_tree_add_48_2_groupi_n_395, csa_tree_add_48_2_groupi_n_396,
     csa_tree_add_48_2_groupi_n_397, csa_tree_add_48_2_groupi_n_398,
     csa_tree_add_48_2_groupi_n_399, csa_tree_add_48_2_groupi_n_400,
     csa_tree_add_48_2_groupi_n_401, csa_tree_add_48_2_groupi_n_402,
     csa_tree_add_48_2_groupi_n_403, csa_tree_add_48_2_groupi_n_404,
     csa_tree_add_48_2_groupi_n_405, csa_tree_add_48_2_groupi_n_406,
     csa_tree_add_48_2_groupi_n_407, csa_tree_add_48_2_groupi_n_408,
     csa_tree_add_48_2_groupi_n_409, csa_tree_add_48_2_groupi_n_410,
     csa_tree_add_48_2_groupi_n_411, csa_tree_add_48_2_groupi_n_412,
     csa_tree_add_48_2_groupi_n_413, csa_tree_add_48_2_groupi_n_414,
     csa_tree_add_48_2_groupi_n_415, csa_tree_add_48_2_groupi_n_416,
     csa_tree_add_48_2_groupi_n_418, csa_tree_add_48_2_groupi_n_419,
     csa_tree_add_48_2_groupi_n_420, csa_tree_add_48_2_groupi_n_421,
     csa_tree_add_48_2_groupi_n_422, csa_tree_add_48_2_groupi_n_423,
     csa_tree_add_48_2_groupi_n_424, csa_tree_add_48_2_groupi_n_425,
     csa_tree_add_48_2_groupi_n_426, csa_tree_add_48_2_groupi_n_427,
     csa_tree_add_48_2_groupi_n_428, csa_tree_add_48_2_groupi_n_430,
     csa_tree_add_48_2_groupi_n_431, csa_tree_add_48_2_groupi_n_432,
     csa_tree_add_48_2_groupi_n_433, csa_tree_add_48_2_groupi_n_434,
     csa_tree_add_48_2_groupi_n_435, csa_tree_add_48_2_groupi_n_436,
     csa_tree_add_48_2_groupi_n_438, csa_tree_add_48_2_groupi_n_439,
     csa_tree_add_48_2_groupi_n_440, csa_tree_add_48_2_groupi_n_441,
     csa_tree_add_48_2_groupi_n_442, csa_tree_add_48_2_groupi_n_443,
     csa_tree_add_48_2_groupi_n_444, csa_tree_add_48_2_groupi_n_445,
     csa_tree_add_48_2_groupi_n_446, csa_tree_add_48_2_groupi_n_447,
     csa_tree_add_48_2_groupi_n_448, csa_tree_add_48_2_groupi_n_449,
     csa_tree_add_48_2_groupi_n_450, csa_tree_add_48_2_groupi_n_451,
     csa_tree_add_48_2_groupi_n_452, csa_tree_add_48_2_groupi_n_453,
     csa_tree_add_48_2_groupi_n_454, csa_tree_add_48_2_groupi_n_455,
     csa_tree_add_48_2_groupi_n_456, csa_tree_add_48_2_groupi_n_457,
     csa_tree_add_48_2_groupi_n_458, csa_tree_add_48_2_groupi_n_459,
     csa_tree_add_48_2_groupi_n_460, csa_tree_add_48_2_groupi_n_461,
     csa_tree_add_48_2_groupi_n_462, csa_tree_add_48_2_groupi_n_463,
     csa_tree_add_48_2_groupi_n_464, csa_tree_add_48_2_groupi_n_465,
     csa_tree_add_48_2_groupi_n_466, csa_tree_add_48_2_groupi_n_467,
     csa_tree_add_48_2_groupi_n_468, csa_tree_add_48_2_groupi_n_469,
     csa_tree_add_48_2_groupi_n_470, csa_tree_add_48_2_groupi_n_471,
     csa_tree_add_48_2_groupi_n_472, csa_tree_add_48_2_groupi_n_473,
     csa_tree_add_48_2_groupi_n_474, csa_tree_add_48_2_groupi_n_475,
     csa_tree_add_48_2_groupi_n_476, csa_tree_add_48_2_groupi_n_477,
     csa_tree_add_48_2_groupi_n_478, csa_tree_add_48_2_groupi_n_479,
     csa_tree_add_48_2_groupi_n_480, csa_tree_add_48_2_groupi_n_481,
     csa_tree_add_48_2_groupi_n_482, csa_tree_add_48_2_groupi_n_483,
     csa_tree_add_48_2_groupi_n_484, csa_tree_add_48_2_groupi_n_485,
     csa_tree_add_48_2_groupi_n_486, csa_tree_add_48_2_groupi_n_487,
     csa_tree_add_48_2_groupi_n_488, csa_tree_add_48_2_groupi_n_489,
     csa_tree_add_48_2_groupi_n_490, csa_tree_add_48_2_groupi_n_491,
     csa_tree_add_48_2_groupi_n_492, csa_tree_add_48_2_groupi_n_493,
     csa_tree_add_48_2_groupi_n_494, csa_tree_add_48_2_groupi_n_495,
     csa_tree_add_48_2_groupi_n_496, csa_tree_add_48_2_groupi_n_497,
     csa_tree_add_48_2_groupi_n_498, csa_tree_add_48_2_groupi_n_499,
     csa_tree_add_48_2_groupi_n_500, csa_tree_add_48_2_groupi_n_501,
     csa_tree_add_48_2_groupi_n_502, csa_tree_add_48_2_groupi_n_503,
     csa_tree_add_48_2_groupi_n_504, csa_tree_add_48_2_groupi_n_505,
     csa_tree_add_48_2_groupi_n_506, csa_tree_add_48_2_groupi_n_507,
     csa_tree_add_48_2_groupi_n_508, csa_tree_add_48_2_groupi_n_509,
     csa_tree_add_48_2_groupi_n_510, csa_tree_add_48_2_groupi_n_511,
     csa_tree_add_48_2_groupi_n_512, csa_tree_add_48_2_groupi_n_513,
     csa_tree_add_48_2_groupi_n_514, csa_tree_add_48_2_groupi_n_515,
     csa_tree_add_48_2_groupi_n_516, csa_tree_add_48_2_groupi_n_517,
     csa_tree_add_48_2_groupi_n_518, csa_tree_add_48_2_groupi_n_519,
     csa_tree_add_48_2_groupi_n_520, csa_tree_add_48_2_groupi_n_521,
     csa_tree_add_48_2_groupi_n_522, csa_tree_add_48_2_groupi_n_523,
     csa_tree_add_48_2_groupi_n_524, csa_tree_add_48_2_groupi_n_525,
     csa_tree_add_48_2_groupi_n_526, csa_tree_add_48_2_groupi_n_527,
     csa_tree_add_48_2_groupi_n_528, csa_tree_add_48_2_groupi_n_529,
     csa_tree_add_48_2_groupi_n_530, csa_tree_add_48_2_groupi_n_531,
     csa_tree_add_48_2_groupi_n_532, csa_tree_add_48_2_groupi_n_533,
     csa_tree_add_48_2_groupi_n_534, csa_tree_add_48_2_groupi_n_535,
     csa_tree_add_48_2_groupi_n_536, csa_tree_add_48_2_groupi_n_537,
     csa_tree_add_48_2_groupi_n_538, csa_tree_add_48_2_groupi_n_539,
     csa_tree_add_48_2_groupi_n_540, csa_tree_add_48_2_groupi_n_541,
     csa_tree_add_48_2_groupi_n_542, csa_tree_add_48_2_groupi_n_543,
     csa_tree_add_48_2_groupi_n_544, csa_tree_add_48_2_groupi_n_545,
     csa_tree_add_48_2_groupi_n_546, csa_tree_add_48_2_groupi_n_547,
     csa_tree_add_48_2_groupi_n_548, csa_tree_add_48_2_groupi_n_549,
     csa_tree_add_48_2_groupi_n_550, csa_tree_add_48_2_groupi_n_551,
     csa_tree_add_48_2_groupi_n_552, csa_tree_add_48_2_groupi_n_553,
     csa_tree_add_48_2_groupi_n_554, csa_tree_add_48_2_groupi_n_555,
     csa_tree_add_48_2_groupi_n_556, csa_tree_add_48_2_groupi_n_557,
     csa_tree_add_48_2_groupi_n_558, csa_tree_add_48_2_groupi_n_559,
     csa_tree_add_48_2_groupi_n_560, csa_tree_add_48_2_groupi_n_561,
     csa_tree_add_48_2_groupi_n_562, csa_tree_add_48_2_groupi_n_563,
     csa_tree_add_48_2_groupi_n_564, csa_tree_add_48_2_groupi_n_565,
     csa_tree_add_48_2_groupi_n_566, csa_tree_add_48_2_groupi_n_567,
     csa_tree_add_48_2_groupi_n_568, csa_tree_add_48_2_groupi_n_569,
     csa_tree_add_48_2_groupi_n_570, csa_tree_add_48_2_groupi_n_571,
     csa_tree_add_48_2_groupi_n_572, csa_tree_add_48_2_groupi_n_573,
     csa_tree_add_48_2_groupi_n_574, csa_tree_add_48_2_groupi_n_575,
     csa_tree_add_48_2_groupi_n_576, csa_tree_add_48_2_groupi_n_577,
     csa_tree_add_48_2_groupi_n_578, csa_tree_add_48_2_groupi_n_579,
     csa_tree_add_48_2_groupi_n_580, csa_tree_add_48_2_groupi_n_581,
     csa_tree_add_48_2_groupi_n_582, csa_tree_add_48_2_groupi_n_583,
     csa_tree_add_48_2_groupi_n_584, csa_tree_add_48_2_groupi_n_585,
     csa_tree_add_48_2_groupi_n_586, csa_tree_add_48_2_groupi_n_587,
     csa_tree_add_48_2_groupi_n_588, csa_tree_add_48_2_groupi_n_589,
     csa_tree_add_48_2_groupi_n_590, csa_tree_add_48_2_groupi_n_591,
     csa_tree_add_48_2_groupi_n_592, csa_tree_add_48_2_groupi_n_593,
     csa_tree_add_48_2_groupi_n_594, csa_tree_add_48_2_groupi_n_595,
     csa_tree_add_48_2_groupi_n_596, csa_tree_add_48_2_groupi_n_597,
     csa_tree_add_48_2_groupi_n_598, csa_tree_add_48_2_groupi_n_599,
     csa_tree_add_48_2_groupi_n_600, csa_tree_add_48_2_groupi_n_601,
     csa_tree_add_48_2_groupi_n_602, csa_tree_add_48_2_groupi_n_603,
     csa_tree_add_48_2_groupi_n_604, csa_tree_add_48_2_groupi_n_605,
     csa_tree_add_48_2_groupi_n_606, csa_tree_add_48_2_groupi_n_607,
     csa_tree_add_48_2_groupi_n_608, csa_tree_add_48_2_groupi_n_609,
     csa_tree_add_48_2_groupi_n_610, csa_tree_add_48_2_groupi_n_611,
     csa_tree_add_48_2_groupi_n_612, csa_tree_add_48_2_groupi_n_613,
     csa_tree_add_48_2_groupi_n_614, csa_tree_add_48_2_groupi_n_615,
     csa_tree_add_48_2_groupi_n_616, csa_tree_add_48_2_groupi_n_617,
     csa_tree_add_48_2_groupi_n_618, csa_tree_add_48_2_groupi_n_619,
     csa_tree_add_48_2_groupi_n_620, csa_tree_add_48_2_groupi_n_621,
     csa_tree_add_48_2_groupi_n_622, csa_tree_add_48_2_groupi_n_623,
     csa_tree_add_48_2_groupi_n_624, csa_tree_add_48_2_groupi_n_625,
     csa_tree_add_48_2_groupi_n_626, csa_tree_add_48_2_groupi_n_627,
     csa_tree_add_48_2_groupi_n_628, csa_tree_add_48_2_groupi_n_629,
     csa_tree_add_48_2_groupi_n_630, csa_tree_add_48_2_groupi_n_631,
     csa_tree_add_48_2_groupi_n_632, csa_tree_add_48_2_groupi_n_633,
     csa_tree_add_48_2_groupi_n_634, csa_tree_add_48_2_groupi_n_635,
     csa_tree_add_48_2_groupi_n_636, csa_tree_add_48_2_groupi_n_637,
     csa_tree_add_48_2_groupi_n_638, csa_tree_add_48_2_groupi_n_639,
     csa_tree_add_48_2_groupi_n_640, csa_tree_add_48_2_groupi_n_641,
     csa_tree_add_48_2_groupi_n_642, csa_tree_add_48_2_groupi_n_643,
     csa_tree_add_48_2_groupi_n_644, csa_tree_add_48_2_groupi_n_645,
     csa_tree_add_48_2_groupi_n_646, csa_tree_add_48_2_groupi_n_647,
     csa_tree_add_48_2_groupi_n_648, csa_tree_add_48_2_groupi_n_649,
     csa_tree_add_48_2_groupi_n_650, csa_tree_add_48_2_groupi_n_651,
     csa_tree_add_48_2_groupi_n_652, csa_tree_add_48_2_groupi_n_653,
     csa_tree_add_48_2_groupi_n_654, csa_tree_add_48_2_groupi_n_655,
     csa_tree_add_48_2_groupi_n_656, csa_tree_add_48_2_groupi_n_657,
     csa_tree_add_48_2_groupi_n_658, csa_tree_add_48_2_groupi_n_659,
     csa_tree_add_48_2_groupi_n_660, csa_tree_add_48_2_groupi_n_661,
     csa_tree_add_48_2_groupi_n_662, csa_tree_add_48_2_groupi_n_663,
     csa_tree_add_48_2_groupi_n_664, csa_tree_add_48_2_groupi_n_665,
     csa_tree_add_48_2_groupi_n_666, csa_tree_add_48_2_groupi_n_667,
     csa_tree_add_48_2_groupi_n_668, csa_tree_add_48_2_groupi_n_669,
     csa_tree_add_48_2_groupi_n_670, csa_tree_add_48_2_groupi_n_671,
     csa_tree_add_48_2_groupi_n_672, csa_tree_add_48_2_groupi_n_673,
     csa_tree_add_48_2_groupi_n_674, csa_tree_add_48_2_groupi_n_675,
     csa_tree_add_48_2_groupi_n_676, csa_tree_add_48_2_groupi_n_677,
     csa_tree_add_48_2_groupi_n_678, csa_tree_add_48_2_groupi_n_679,
     csa_tree_add_48_2_groupi_n_680, csa_tree_add_48_2_groupi_n_681,
     csa_tree_add_48_2_groupi_n_682, csa_tree_add_48_2_groupi_n_683,
     csa_tree_add_48_2_groupi_n_684, csa_tree_add_48_2_groupi_n_685,
     csa_tree_add_48_2_groupi_n_686, csa_tree_add_48_2_groupi_n_687,
     csa_tree_add_48_2_groupi_n_688, csa_tree_add_48_2_groupi_n_689,
     csa_tree_add_48_2_groupi_n_690, csa_tree_add_48_2_groupi_n_691,
     csa_tree_add_48_2_groupi_n_692, csa_tree_add_48_2_groupi_n_693,
     csa_tree_add_48_2_groupi_n_694, csa_tree_add_48_2_groupi_n_695,
     csa_tree_add_48_2_groupi_n_696, csa_tree_add_48_2_groupi_n_697,
     csa_tree_add_48_2_groupi_n_698, csa_tree_add_48_2_groupi_n_699,
     csa_tree_add_48_2_groupi_n_700, csa_tree_add_48_2_groupi_n_701,
     csa_tree_add_48_2_groupi_n_702, csa_tree_add_48_2_groupi_n_703,
     csa_tree_add_48_2_groupi_n_704, csa_tree_add_48_2_groupi_n_705,
     csa_tree_add_48_2_groupi_n_706, csa_tree_add_48_2_groupi_n_707,
     csa_tree_add_48_2_groupi_n_708, csa_tree_add_48_2_groupi_n_709,
     csa_tree_add_48_2_groupi_n_710, csa_tree_add_48_2_groupi_n_711,
     csa_tree_add_48_2_groupi_n_712, csa_tree_add_48_2_groupi_n_713,
     csa_tree_add_48_2_groupi_n_714, csa_tree_add_48_2_groupi_n_715,
     csa_tree_add_48_2_groupi_n_716, csa_tree_add_48_2_groupi_n_717,
     csa_tree_add_48_2_groupi_n_718, csa_tree_add_48_2_groupi_n_719,
     csa_tree_add_48_2_groupi_n_720, csa_tree_add_48_2_groupi_n_721,
     csa_tree_add_48_2_groupi_n_722, csa_tree_add_48_2_groupi_n_723,
     csa_tree_add_48_2_groupi_n_724, csa_tree_add_48_2_groupi_n_725,
     csa_tree_add_48_2_groupi_n_726, csa_tree_add_48_2_groupi_n_727,
     csa_tree_add_48_2_groupi_n_728, csa_tree_add_48_2_groupi_n_729,
     csa_tree_add_48_2_groupi_n_730, csa_tree_add_48_2_groupi_n_731,
     csa_tree_add_48_2_groupi_n_732, csa_tree_add_48_2_groupi_n_733,
     csa_tree_add_48_2_groupi_n_734, csa_tree_add_48_2_groupi_n_735,
     csa_tree_add_48_2_groupi_n_736, csa_tree_add_48_2_groupi_n_737,
     csa_tree_add_48_2_groupi_n_738, csa_tree_add_48_2_groupi_n_739,
     csa_tree_add_48_2_groupi_n_740, csa_tree_add_48_2_groupi_n_741,
     csa_tree_add_48_2_groupi_n_742, csa_tree_add_48_2_groupi_n_743,
     csa_tree_add_48_2_groupi_n_744, csa_tree_add_48_2_groupi_n_745,
     csa_tree_add_48_2_groupi_n_746, csa_tree_add_48_2_groupi_n_747,
     csa_tree_add_48_2_groupi_n_748, csa_tree_add_48_2_groupi_n_749,
     csa_tree_add_48_2_groupi_n_750, csa_tree_add_48_2_groupi_n_751,
     csa_tree_add_48_2_groupi_n_752, csa_tree_add_48_2_groupi_n_753,
     csa_tree_add_48_2_groupi_n_754, csa_tree_add_48_2_groupi_n_755,
     csa_tree_add_48_2_groupi_n_756, csa_tree_add_48_2_groupi_n_757,
     csa_tree_add_48_2_groupi_n_758, csa_tree_add_48_2_groupi_n_759,
     csa_tree_add_48_2_groupi_n_760, csa_tree_add_48_2_groupi_n_761,
     csa_tree_add_48_2_groupi_n_762, csa_tree_add_48_2_groupi_n_763,
     csa_tree_add_48_2_groupi_n_764, csa_tree_add_48_2_groupi_n_765,
     csa_tree_add_48_2_groupi_n_766, csa_tree_add_48_2_groupi_n_767,
     csa_tree_add_48_2_groupi_n_768, csa_tree_add_48_2_groupi_n_769,
     csa_tree_add_48_2_groupi_n_770, csa_tree_add_48_2_groupi_n_771,
     csa_tree_add_48_2_groupi_n_772, csa_tree_add_48_2_groupi_n_773,
     csa_tree_add_48_2_groupi_n_774, csa_tree_add_48_2_groupi_n_775,
     csa_tree_add_48_2_groupi_n_776, csa_tree_add_48_2_groupi_n_777,
     csa_tree_add_48_2_groupi_n_778, csa_tree_add_48_2_groupi_n_779,
     csa_tree_add_48_2_groupi_n_780, csa_tree_add_48_2_groupi_n_781,
     csa_tree_add_48_2_groupi_n_782, csa_tree_add_48_2_groupi_n_783,
     csa_tree_add_48_2_groupi_n_784, csa_tree_add_48_2_groupi_n_785,
     csa_tree_add_48_2_groupi_n_786, csa_tree_add_48_2_groupi_n_787,
     csa_tree_add_48_2_groupi_n_788, csa_tree_add_48_2_groupi_n_789,
     csa_tree_add_48_2_groupi_n_790, csa_tree_add_48_2_groupi_n_791,
     csa_tree_add_48_2_groupi_n_792, csa_tree_add_48_2_groupi_n_793,
     csa_tree_add_48_2_groupi_n_794, csa_tree_add_48_2_groupi_n_795,
     csa_tree_add_48_2_groupi_n_796, csa_tree_add_48_2_groupi_n_797,
     csa_tree_add_48_2_groupi_n_798, csa_tree_add_48_2_groupi_n_799,
     csa_tree_add_48_2_groupi_n_800, csa_tree_add_48_2_groupi_n_801,
     csa_tree_add_48_2_groupi_n_802, csa_tree_add_48_2_groupi_n_803,
     csa_tree_add_48_2_groupi_n_804, csa_tree_add_48_2_groupi_n_805,
     csa_tree_add_48_2_groupi_n_806, csa_tree_add_48_2_groupi_n_807,
     csa_tree_add_48_2_groupi_n_808, csa_tree_add_48_2_groupi_n_809,
     csa_tree_add_48_2_groupi_n_810, csa_tree_add_48_2_groupi_n_811,
     csa_tree_add_48_2_groupi_n_812, csa_tree_add_48_2_groupi_n_813,
     csa_tree_add_48_2_groupi_n_814, csa_tree_add_48_2_groupi_n_815,
     csa_tree_add_48_2_groupi_n_816, csa_tree_add_48_2_groupi_n_817,
     csa_tree_add_48_2_groupi_n_818, csa_tree_add_48_2_groupi_n_819,
     csa_tree_add_48_2_groupi_n_820, csa_tree_add_48_2_groupi_n_821,
     csa_tree_add_48_2_groupi_n_822, csa_tree_add_48_2_groupi_n_823,
     csa_tree_add_48_2_groupi_n_824, csa_tree_add_48_2_groupi_n_825,
     csa_tree_add_48_2_groupi_n_826, csa_tree_add_48_2_groupi_n_827,
     csa_tree_add_48_2_groupi_n_828, csa_tree_add_48_2_groupi_n_829,
     csa_tree_add_48_2_groupi_n_830, csa_tree_add_48_2_groupi_n_831,
     csa_tree_add_48_2_groupi_n_832, csa_tree_add_48_2_groupi_n_833,
     csa_tree_add_48_2_groupi_n_834, csa_tree_add_48_2_groupi_n_835,
     csa_tree_add_48_2_groupi_n_836, csa_tree_add_48_2_groupi_n_837,
     csa_tree_add_48_2_groupi_n_838, csa_tree_add_48_2_groupi_n_839,
     csa_tree_add_48_2_groupi_n_840, csa_tree_add_48_2_groupi_n_841,
     csa_tree_add_48_2_groupi_n_842, csa_tree_add_48_2_groupi_n_843,
     csa_tree_add_48_2_groupi_n_844, csa_tree_add_48_2_groupi_n_845,
     csa_tree_add_48_2_groupi_n_846, csa_tree_add_48_2_groupi_n_847,
     csa_tree_add_48_2_groupi_n_848, csa_tree_add_48_2_groupi_n_850,
     csa_tree_add_48_2_groupi_n_851, csa_tree_add_48_2_groupi_n_852,
     csa_tree_add_48_2_groupi_n_853, csa_tree_add_48_2_groupi_n_854,
     csa_tree_add_48_2_groupi_n_855, csa_tree_add_48_2_groupi_n_856,
     csa_tree_add_48_2_groupi_n_857, csa_tree_add_48_2_groupi_n_858,
     csa_tree_add_48_2_groupi_n_859, csa_tree_add_48_2_groupi_n_860,
     csa_tree_add_48_2_groupi_n_861, csa_tree_add_48_2_groupi_n_862,
     csa_tree_add_48_2_groupi_n_863, csa_tree_add_48_2_groupi_n_864,
     csa_tree_add_48_2_groupi_n_865, csa_tree_add_48_2_groupi_n_866,
     csa_tree_add_48_2_groupi_n_867, csa_tree_add_48_2_groupi_n_868,
     csa_tree_add_48_2_groupi_n_869, csa_tree_add_48_2_groupi_n_870,
     csa_tree_add_48_2_groupi_n_871, csa_tree_add_48_2_groupi_n_872,
     csa_tree_add_48_2_groupi_n_873, csa_tree_add_48_2_groupi_n_874,
     csa_tree_add_48_2_groupi_n_875, csa_tree_add_48_2_groupi_n_876,
     csa_tree_add_48_2_groupi_n_877, csa_tree_add_48_2_groupi_n_878,
     csa_tree_add_48_2_groupi_n_879, csa_tree_add_48_2_groupi_n_880,
     csa_tree_add_48_2_groupi_n_881, csa_tree_add_48_2_groupi_n_882,
     csa_tree_add_48_2_groupi_n_883, csa_tree_add_48_2_groupi_n_884,
     csa_tree_add_48_2_groupi_n_885, csa_tree_add_48_2_groupi_n_886,
     csa_tree_add_48_2_groupi_n_887, csa_tree_add_48_2_groupi_n_888,
     csa_tree_add_48_2_groupi_n_889, csa_tree_add_48_2_groupi_n_890,
     csa_tree_add_48_2_groupi_n_891, csa_tree_add_48_2_groupi_n_892,
     csa_tree_add_48_2_groupi_n_893, csa_tree_add_48_2_groupi_n_894,
     csa_tree_add_48_2_groupi_n_895, csa_tree_add_48_2_groupi_n_896,
     csa_tree_add_48_2_groupi_n_897, csa_tree_add_48_2_groupi_n_898,
     csa_tree_add_48_2_groupi_n_899, csa_tree_add_48_2_groupi_n_900,
     csa_tree_add_48_2_groupi_n_901, csa_tree_add_48_2_groupi_n_902,
     csa_tree_add_48_2_groupi_n_903, csa_tree_add_48_2_groupi_n_904,
     csa_tree_add_48_2_groupi_n_905, csa_tree_add_48_2_groupi_n_906,
     csa_tree_add_48_2_groupi_n_907, csa_tree_add_48_2_groupi_n_908,
     csa_tree_add_48_2_groupi_n_909, csa_tree_add_48_2_groupi_n_910,
     csa_tree_add_48_2_groupi_n_911, csa_tree_add_48_2_groupi_n_912,
     csa_tree_add_48_2_groupi_n_913, csa_tree_add_48_2_groupi_n_914,
     csa_tree_add_48_2_groupi_n_915, csa_tree_add_48_2_groupi_n_916,
     csa_tree_add_48_2_groupi_n_917, csa_tree_add_48_2_groupi_n_918,
     csa_tree_add_48_2_groupi_n_919, csa_tree_add_48_2_groupi_n_920,
     csa_tree_add_48_2_groupi_n_921, csa_tree_add_48_2_groupi_n_922,
     csa_tree_add_48_2_groupi_n_923, csa_tree_add_48_2_groupi_n_924,
     csa_tree_add_48_2_groupi_n_925, csa_tree_add_48_2_groupi_n_926,
     csa_tree_add_48_2_groupi_n_927, csa_tree_add_48_2_groupi_n_928,
     csa_tree_add_48_2_groupi_n_929, csa_tree_add_48_2_groupi_n_930,
     csa_tree_add_48_2_groupi_n_931, csa_tree_add_48_2_groupi_n_932,
     csa_tree_add_48_2_groupi_n_933, csa_tree_add_48_2_groupi_n_934,
     csa_tree_add_48_2_groupi_n_935, csa_tree_add_48_2_groupi_n_936,
     csa_tree_add_48_2_groupi_n_937, csa_tree_add_48_2_groupi_n_938,
     csa_tree_add_48_2_groupi_n_939, csa_tree_add_48_2_groupi_n_940,
     csa_tree_add_48_2_groupi_n_941, csa_tree_add_48_2_groupi_n_942,
     csa_tree_add_48_2_groupi_n_943, csa_tree_add_48_2_groupi_n_944,
     csa_tree_add_48_2_groupi_n_945, csa_tree_add_48_2_groupi_n_946,
     csa_tree_add_48_2_groupi_n_947, csa_tree_add_48_2_groupi_n_948,
     csa_tree_add_48_2_groupi_n_949, csa_tree_add_48_2_groupi_n_950,
     csa_tree_add_48_2_groupi_n_951, csa_tree_add_48_2_groupi_n_952,
     csa_tree_add_48_2_groupi_n_953, csa_tree_add_48_2_groupi_n_954,
     csa_tree_add_48_2_groupi_n_955, csa_tree_add_48_2_groupi_n_956,
     csa_tree_add_48_2_groupi_n_957, csa_tree_add_48_2_groupi_n_958,
     csa_tree_add_48_2_groupi_n_959, csa_tree_add_48_2_groupi_n_960,
     csa_tree_add_48_2_groupi_n_961, csa_tree_add_48_2_groupi_n_962,
     csa_tree_add_48_2_groupi_n_963, csa_tree_add_48_2_groupi_n_964,
     csa_tree_add_48_2_groupi_n_965, csa_tree_add_48_2_groupi_n_966,
     csa_tree_add_48_2_groupi_n_967, csa_tree_add_48_2_groupi_n_968,
     csa_tree_add_48_2_groupi_n_969, csa_tree_add_48_2_groupi_n_970,
     csa_tree_add_48_2_groupi_n_971, csa_tree_add_48_2_groupi_n_972,
     csa_tree_add_48_2_groupi_n_973, csa_tree_add_48_2_groupi_n_974,
     csa_tree_add_48_2_groupi_n_975, csa_tree_add_48_2_groupi_n_976,
     csa_tree_add_48_2_groupi_n_977, csa_tree_add_48_2_groupi_n_978,
     csa_tree_add_48_2_groupi_n_979, csa_tree_add_48_2_groupi_n_980,
     csa_tree_add_48_2_groupi_n_981, csa_tree_add_48_2_groupi_n_982,
     csa_tree_add_48_2_groupi_n_983, csa_tree_add_48_2_groupi_n_984,
     csa_tree_add_48_2_groupi_n_985, csa_tree_add_48_2_groupi_n_986,
     csa_tree_add_48_2_groupi_n_987, csa_tree_add_48_2_groupi_n_988,
     csa_tree_add_48_2_groupi_n_989, csa_tree_add_48_2_groupi_n_990,
     csa_tree_add_48_2_groupi_n_991, csa_tree_add_48_2_groupi_n_992,
     csa_tree_add_48_2_groupi_n_993, csa_tree_add_48_2_groupi_n_994,
     csa_tree_add_48_2_groupi_n_995, csa_tree_add_48_2_groupi_n_996,
     csa_tree_add_48_2_groupi_n_997, csa_tree_add_48_2_groupi_n_998,
     csa_tree_add_48_2_groupi_n_999, csa_tree_add_48_2_groupi_n_1000,
     csa_tree_add_48_2_groupi_n_1001, csa_tree_add_48_2_groupi_n_1002,
     csa_tree_add_48_2_groupi_n_1003, csa_tree_add_48_2_groupi_n_1004,
     csa_tree_add_48_2_groupi_n_1005, csa_tree_add_48_2_groupi_n_1006,
     csa_tree_add_48_2_groupi_n_1007, csa_tree_add_48_2_groupi_n_1008,
     csa_tree_add_48_2_groupi_n_1009, csa_tree_add_48_2_groupi_n_1010,
     csa_tree_add_48_2_groupi_n_1011, csa_tree_add_48_2_groupi_n_1012,
     csa_tree_add_48_2_groupi_n_1013, csa_tree_add_48_2_groupi_n_1014,
     csa_tree_add_48_2_groupi_n_1015, csa_tree_add_48_2_groupi_n_1016,
     csa_tree_add_48_2_groupi_n_1017, csa_tree_add_48_2_groupi_n_1018,
     csa_tree_add_48_2_groupi_n_1019, csa_tree_add_48_2_groupi_n_1020,
     csa_tree_add_48_2_groupi_n_1021, csa_tree_add_48_2_groupi_n_1022,
     csa_tree_add_48_2_groupi_n_1023, csa_tree_add_48_2_groupi_n_1024,
     csa_tree_add_48_2_groupi_n_1025, csa_tree_add_48_2_groupi_n_1026,
     csa_tree_add_48_2_groupi_n_1027, csa_tree_add_48_2_groupi_n_1028,
     csa_tree_add_48_2_groupi_n_1029, csa_tree_add_48_2_groupi_n_1030,
     csa_tree_add_48_2_groupi_n_1031, csa_tree_add_48_2_groupi_n_1032,
     csa_tree_add_48_2_groupi_n_1033, csa_tree_add_48_2_groupi_n_1034,
     csa_tree_add_48_2_groupi_n_1035, csa_tree_add_48_2_groupi_n_1036,
     csa_tree_add_48_2_groupi_n_1037, csa_tree_add_48_2_groupi_n_1038,
     csa_tree_add_48_2_groupi_n_1039, csa_tree_add_48_2_groupi_n_1040,
     csa_tree_add_48_2_groupi_n_1041, csa_tree_add_48_2_groupi_n_1042,
     csa_tree_add_48_2_groupi_n_1043, csa_tree_add_48_2_groupi_n_1044,
     csa_tree_add_48_2_groupi_n_1045, csa_tree_add_48_2_groupi_n_1046,
     csa_tree_add_48_2_groupi_n_1047, csa_tree_add_48_2_groupi_n_1048,
     csa_tree_add_48_2_groupi_n_1049, csa_tree_add_48_2_groupi_n_1050,
     csa_tree_add_48_2_groupi_n_1052, csa_tree_add_48_2_groupi_n_1053,
     csa_tree_add_48_2_groupi_n_1054, csa_tree_add_48_2_groupi_n_1055,
     csa_tree_add_48_2_groupi_n_1056, csa_tree_add_48_2_groupi_n_1057,
     csa_tree_add_48_2_groupi_n_1058, csa_tree_add_48_2_groupi_n_1059,
     csa_tree_add_48_2_groupi_n_1060, csa_tree_add_48_2_groupi_n_1061,
     csa_tree_add_48_2_groupi_n_1062, csa_tree_add_48_2_groupi_n_1063,
     csa_tree_add_48_2_groupi_n_1064, csa_tree_add_48_2_groupi_n_1066,
     csa_tree_add_48_2_groupi_n_1067, csa_tree_add_48_2_groupi_n_1070,
     csa_tree_add_48_2_groupi_n_1071, csa_tree_add_48_2_groupi_n_1072,
     csa_tree_add_48_2_groupi_n_1073, csa_tree_add_48_2_groupi_n_1074,
     csa_tree_add_48_2_groupi_n_1075, csa_tree_add_48_2_groupi_n_1076,
     csa_tree_add_48_2_groupi_n_1077, csa_tree_add_48_2_groupi_n_1078,
     csa_tree_add_48_2_groupi_n_1079, csa_tree_add_48_2_groupi_n_1080,
     csa_tree_add_48_2_groupi_n_1081, csa_tree_add_48_2_groupi_n_1082,
     csa_tree_add_48_2_groupi_n_1083, csa_tree_add_48_2_groupi_n_1084,
     csa_tree_add_48_2_groupi_n_1085, csa_tree_add_48_2_groupi_n_1086,
     csa_tree_add_48_2_groupi_n_1087, csa_tree_add_48_2_groupi_n_1088,
     csa_tree_add_48_2_groupi_n_1089, csa_tree_add_48_2_groupi_n_1090,
     csa_tree_add_48_2_groupi_n_1091, csa_tree_add_48_2_groupi_n_1092,
     csa_tree_add_48_2_groupi_n_1093, csa_tree_add_48_2_groupi_n_1094,
     csa_tree_add_48_2_groupi_n_1095, csa_tree_add_48_2_groupi_n_1096,
     csa_tree_add_48_2_groupi_n_1097, csa_tree_add_48_2_groupi_n_1099,
     csa_tree_add_48_2_groupi_n_1100, csa_tree_add_48_2_groupi_n_1101,
     csa_tree_add_48_2_groupi_n_1102, csa_tree_add_48_2_groupi_n_1103,
     csa_tree_add_48_2_groupi_n_1104, csa_tree_add_48_2_groupi_n_1105,
     csa_tree_add_48_2_groupi_n_1106, csa_tree_add_48_2_groupi_n_1107,
     csa_tree_add_48_2_groupi_n_1109, csa_tree_add_48_2_groupi_n_1110,
     csa_tree_add_48_2_groupi_n_1111, csa_tree_add_48_2_groupi_n_1112,
     csa_tree_add_48_2_groupi_n_1113, csa_tree_add_48_2_groupi_n_1114,
     csa_tree_add_48_2_groupi_n_1115, csa_tree_add_48_2_groupi_n_1116,
     csa_tree_add_48_2_groupi_n_1117, csa_tree_add_48_2_groupi_n_1118,
     csa_tree_add_48_2_groupi_n_1119, csa_tree_add_48_2_groupi_n_1120,
     csa_tree_add_48_2_groupi_n_1121, csa_tree_add_48_2_groupi_n_1122,
     csa_tree_add_48_2_groupi_n_1124, csa_tree_add_48_2_groupi_n_1125,
     csa_tree_add_48_2_groupi_n_1126, csa_tree_add_48_2_groupi_n_1127,
     csa_tree_add_48_2_groupi_n_1128, csa_tree_add_48_2_groupi_n_1129,
     csa_tree_add_48_2_groupi_n_1130, csa_tree_add_48_2_groupi_n_1131,
     csa_tree_add_48_2_groupi_n_1132, csa_tree_add_48_2_groupi_n_1133,
     csa_tree_add_48_2_groupi_n_1135, csa_tree_add_48_2_groupi_n_1136,
     csa_tree_add_48_2_groupi_n_1137, csa_tree_add_48_2_groupi_n_1138,
     csa_tree_add_48_2_groupi_n_1139, csa_tree_add_48_2_groupi_n_1140,
     csa_tree_add_48_2_groupi_n_1141, csa_tree_add_48_2_groupi_n_1142,
     csa_tree_add_48_2_groupi_n_1143, csa_tree_add_48_2_groupi_n_1144,
     csa_tree_add_48_2_groupi_n_1145, csa_tree_add_48_2_groupi_n_1146,
     csa_tree_add_48_2_groupi_n_1147, csa_tree_add_48_2_groupi_n_1148,
     csa_tree_add_48_2_groupi_n_1149, csa_tree_add_48_2_groupi_n_1150,
     csa_tree_add_48_2_groupi_n_1151, csa_tree_add_48_2_groupi_n_1152,
     csa_tree_add_48_2_groupi_n_1153, csa_tree_add_48_2_groupi_n_1154,
     csa_tree_add_48_2_groupi_n_1155, csa_tree_add_48_2_groupi_n_1156,
     csa_tree_add_48_2_groupi_n_1157, csa_tree_add_48_2_groupi_n_1158,
     csa_tree_add_48_2_groupi_n_1159, csa_tree_add_48_2_groupi_n_1160,
     csa_tree_add_48_2_groupi_n_1161, csa_tree_add_48_2_groupi_n_1162,
     csa_tree_add_48_2_groupi_n_1163, csa_tree_add_48_2_groupi_n_1164,
     csa_tree_add_48_2_groupi_n_1165, csa_tree_add_48_2_groupi_n_1166,
     csa_tree_add_48_2_groupi_n_1167, csa_tree_add_48_2_groupi_n_1168,
     csa_tree_add_48_2_groupi_n_1169, csa_tree_add_48_2_groupi_n_1170,
     csa_tree_add_48_2_groupi_n_1171, csa_tree_add_48_2_groupi_n_1172,
     csa_tree_add_48_2_groupi_n_1173, csa_tree_add_48_2_groupi_n_1174,
     csa_tree_add_48_2_groupi_n_1175, csa_tree_add_48_2_groupi_n_1176,
     csa_tree_add_48_2_groupi_n_1177, csa_tree_add_48_2_groupi_n_1178,
     csa_tree_add_48_2_groupi_n_1179, csa_tree_add_48_2_groupi_n_1180,
     csa_tree_add_48_2_groupi_n_1181, csa_tree_add_48_2_groupi_n_1182,
     csa_tree_add_48_2_groupi_n_1183, csa_tree_add_48_2_groupi_n_1184,
     csa_tree_add_48_2_groupi_n_1185, csa_tree_add_48_2_groupi_n_1186,
     csa_tree_add_48_2_groupi_n_1189, csa_tree_add_48_2_groupi_n_1190,
     csa_tree_add_48_2_groupi_n_1191, csa_tree_add_48_2_groupi_n_1192,
     csa_tree_add_48_2_groupi_n_1193, csa_tree_add_48_2_groupi_n_1194,
     csa_tree_add_48_2_groupi_n_1195, csa_tree_add_48_2_groupi_n_1196,
     csa_tree_add_48_2_groupi_n_1197, csa_tree_add_48_2_groupi_n_1198,
     csa_tree_add_48_2_groupi_n_1199, csa_tree_add_48_2_groupi_n_1200,
     csa_tree_add_48_2_groupi_n_1201, csa_tree_add_48_2_groupi_n_1202,
     csa_tree_add_48_2_groupi_n_1203, csa_tree_add_48_2_groupi_n_1204,
     csa_tree_add_48_2_groupi_n_1205, csa_tree_add_48_2_groupi_n_1206,
     csa_tree_add_48_2_groupi_n_1207, csa_tree_add_48_2_groupi_n_1208,
     csa_tree_add_48_2_groupi_n_1209, csa_tree_add_48_2_groupi_n_1210,
     csa_tree_add_48_2_groupi_n_1211, csa_tree_add_48_2_groupi_n_1212,
     csa_tree_add_48_2_groupi_n_1213, csa_tree_add_48_2_groupi_n_1214,
     csa_tree_add_48_2_groupi_n_1215, csa_tree_add_48_2_groupi_n_1216,
     csa_tree_add_48_2_groupi_n_1217, csa_tree_add_48_2_groupi_n_1218,
     csa_tree_add_48_2_groupi_n_1219, csa_tree_add_48_2_groupi_n_1220,
     csa_tree_add_48_2_groupi_n_1221, csa_tree_add_48_2_groupi_n_1222,
     csa_tree_add_48_2_groupi_n_1223, csa_tree_add_48_2_groupi_n_1224,
     csa_tree_add_48_2_groupi_n_1225, csa_tree_add_48_2_groupi_n_1226,
     csa_tree_add_48_2_groupi_n_1227, csa_tree_add_48_2_groupi_n_1228,
     csa_tree_add_48_2_groupi_n_1229, csa_tree_add_48_2_groupi_n_1230,
     csa_tree_add_48_2_groupi_n_1231, csa_tree_add_48_2_groupi_n_1232,
     csa_tree_add_48_2_groupi_n_1233, csa_tree_add_48_2_groupi_n_1234,
     csa_tree_add_48_2_groupi_n_1235, csa_tree_add_48_2_groupi_n_1236,
     csa_tree_add_48_2_groupi_n_1237, csa_tree_add_48_2_groupi_n_1238,
     csa_tree_add_48_2_groupi_n_1239, csa_tree_add_48_2_groupi_n_1240,
     csa_tree_add_48_2_groupi_n_1241, csa_tree_add_48_2_groupi_n_1242,
     csa_tree_add_48_2_groupi_n_1243, csa_tree_add_48_2_groupi_n_1244,
     csa_tree_add_48_2_groupi_n_1245, csa_tree_add_48_2_groupi_n_1246,
     csa_tree_add_48_2_groupi_n_1247, csa_tree_add_48_2_groupi_n_1248,
     csa_tree_add_48_2_groupi_n_1249, csa_tree_add_48_2_groupi_n_1250,
     csa_tree_add_48_2_groupi_n_1251, csa_tree_add_48_2_groupi_n_1252,
     csa_tree_add_48_2_groupi_n_1253, csa_tree_add_48_2_groupi_n_1254,
     csa_tree_add_48_2_groupi_n_1255, csa_tree_add_48_2_groupi_n_1256,
     csa_tree_add_48_2_groupi_n_1257, csa_tree_add_48_2_groupi_n_1258,
     csa_tree_add_48_2_groupi_n_1259, csa_tree_add_48_2_groupi_n_1260,
     csa_tree_add_48_2_groupi_n_1261, csa_tree_add_48_2_groupi_n_1262,
     csa_tree_add_48_2_groupi_n_1263, csa_tree_add_48_2_groupi_n_1264,
     csa_tree_add_48_2_groupi_n_1265, csa_tree_add_48_2_groupi_n_1266,
     csa_tree_add_48_2_groupi_n_1267, csa_tree_add_48_2_groupi_n_1268,
     csa_tree_add_48_2_groupi_n_1270, csa_tree_add_48_2_groupi_n_1271,
     csa_tree_add_48_2_groupi_n_1272, csa_tree_add_48_2_groupi_n_1273,
     csa_tree_add_48_2_groupi_n_1274, csa_tree_add_48_2_groupi_n_1275,
     csa_tree_add_48_2_groupi_n_1276, csa_tree_add_48_2_groupi_n_1277,
     csa_tree_add_48_2_groupi_n_1278, csa_tree_add_48_2_groupi_n_1280,
     csa_tree_add_48_2_groupi_n_1281, csa_tree_add_48_2_groupi_n_1282,
     csa_tree_add_48_2_groupi_n_1283, csa_tree_add_48_2_groupi_n_1284,
     csa_tree_add_48_2_groupi_n_1285, csa_tree_add_48_2_groupi_n_1286,
     csa_tree_add_48_2_groupi_n_1287, csa_tree_add_48_2_groupi_n_1288,
     csa_tree_add_48_2_groupi_n_1289, csa_tree_add_48_2_groupi_n_1290,
     csa_tree_add_48_2_groupi_n_1291, csa_tree_add_48_2_groupi_n_1292,
     csa_tree_add_48_2_groupi_n_1293, csa_tree_add_48_2_groupi_n_1294,
     csa_tree_add_48_2_groupi_n_1295, csa_tree_add_48_2_groupi_n_1296,
     csa_tree_add_48_2_groupi_n_1297, csa_tree_add_48_2_groupi_n_1298,
     csa_tree_add_48_2_groupi_n_1299, csa_tree_add_48_2_groupi_n_1300,
     csa_tree_add_48_2_groupi_n_1301, csa_tree_add_48_2_groupi_n_1302,
     csa_tree_add_48_2_groupi_n_1303, csa_tree_add_48_2_groupi_n_1304,
     csa_tree_add_48_2_groupi_n_1305, csa_tree_add_48_2_groupi_n_1307,
     csa_tree_add_48_2_groupi_n_1308, csa_tree_add_48_2_groupi_n_1309,
     csa_tree_add_48_2_groupi_n_1310, csa_tree_add_48_2_groupi_n_1311,
     csa_tree_add_48_2_groupi_n_1312, csa_tree_add_48_2_groupi_n_1313,
     csa_tree_add_48_2_groupi_n_1314, csa_tree_add_48_2_groupi_n_1315,
     csa_tree_add_48_2_groupi_n_1316, csa_tree_add_48_2_groupi_n_1317,
     csa_tree_add_48_2_groupi_n_1318, csa_tree_add_48_2_groupi_n_1319,
     csa_tree_add_48_2_groupi_n_1320, csa_tree_add_48_2_groupi_n_1321,
     csa_tree_add_48_2_groupi_n_1322, csa_tree_add_48_2_groupi_n_1323,
     csa_tree_add_48_2_groupi_n_1324, csa_tree_add_48_2_groupi_n_1325,
     csa_tree_add_48_2_groupi_n_1326, csa_tree_add_48_2_groupi_n_1328,
     csa_tree_add_48_2_groupi_n_1329, csa_tree_add_48_2_groupi_n_1330,
     csa_tree_add_48_2_groupi_n_1331, csa_tree_add_48_2_groupi_n_1332,
     csa_tree_add_48_2_groupi_n_1333, csa_tree_add_48_2_groupi_n_1334,
     csa_tree_add_48_2_groupi_n_1335, csa_tree_add_48_2_groupi_n_1336,
     csa_tree_add_48_2_groupi_n_1337, csa_tree_add_48_2_groupi_n_1338,
     csa_tree_add_48_2_groupi_n_1339, csa_tree_add_48_2_groupi_n_1340,
     csa_tree_add_48_2_groupi_n_1341, csa_tree_add_48_2_groupi_n_1345,
     csa_tree_add_48_2_groupi_n_1346, csa_tree_add_48_2_groupi_n_1347,
     csa_tree_add_48_2_groupi_n_1348, csa_tree_add_48_2_groupi_n_1349,
     csa_tree_add_48_2_groupi_n_1350, csa_tree_add_48_2_groupi_n_1351,
     csa_tree_add_48_2_groupi_n_1352, csa_tree_add_48_2_groupi_n_1353,
     csa_tree_add_48_2_groupi_n_1354, csa_tree_add_48_2_groupi_n_1355,
     csa_tree_add_48_2_groupi_n_1356, csa_tree_add_48_2_groupi_n_1357,
     csa_tree_add_48_2_groupi_n_1358, csa_tree_add_48_2_groupi_n_1359,
     csa_tree_add_48_2_groupi_n_1360, csa_tree_add_48_2_groupi_n_1361,
     csa_tree_add_48_2_groupi_n_1363, csa_tree_add_48_2_groupi_n_1364,
     csa_tree_add_48_2_groupi_n_1365, csa_tree_add_48_2_groupi_n_1366,
     csa_tree_add_48_2_groupi_n_1367, csa_tree_add_48_2_groupi_n_1368,
     csa_tree_add_48_2_groupi_n_1370, csa_tree_add_48_2_groupi_n_1371,
     csa_tree_add_48_2_groupi_n_1372, csa_tree_add_48_2_groupi_n_1373,
     csa_tree_add_48_2_groupi_n_1374, csa_tree_add_48_2_groupi_n_1375,
     csa_tree_add_48_2_groupi_n_1376, csa_tree_add_48_2_groupi_n_1377,
     csa_tree_add_48_2_groupi_n_1378, csa_tree_add_48_2_groupi_n_1379,
     csa_tree_add_48_2_groupi_n_1380, csa_tree_add_48_2_groupi_n_1381,
     csa_tree_add_48_2_groupi_n_1382, csa_tree_add_48_2_groupi_n_1383,
     csa_tree_add_48_2_groupi_n_1384, csa_tree_add_48_2_groupi_n_1386,
     csa_tree_add_48_2_groupi_n_1387, csa_tree_add_48_2_groupi_n_1388,
     csa_tree_add_48_2_groupi_n_1389, csa_tree_add_48_2_groupi_n_1390,
     csa_tree_add_48_2_groupi_n_1391, csa_tree_add_48_2_groupi_n_1392,
     csa_tree_add_48_2_groupi_n_1393, csa_tree_add_48_2_groupi_n_1394,
     csa_tree_add_48_2_groupi_n_1395, csa_tree_add_48_2_groupi_n_1396,
     csa_tree_add_48_2_groupi_n_1397, csa_tree_add_48_2_groupi_n_1398,
     csa_tree_add_48_2_groupi_n_1399, csa_tree_add_48_2_groupi_n_1400,
     csa_tree_add_48_2_groupi_n_1401, csa_tree_add_48_2_groupi_n_1402,
     csa_tree_add_48_2_groupi_n_1403, csa_tree_add_48_2_groupi_n_1404,
     csa_tree_add_48_2_groupi_n_1405, csa_tree_add_48_2_groupi_n_1406,
     csa_tree_add_48_2_groupi_n_1407, csa_tree_add_48_2_groupi_n_1408,
     csa_tree_add_48_2_groupi_n_1409, csa_tree_add_48_2_groupi_n_1410,
     csa_tree_add_48_2_groupi_n_1411, csa_tree_add_48_2_groupi_n_1412,
     csa_tree_add_48_2_groupi_n_1413, csa_tree_add_48_2_groupi_n_1414,
     csa_tree_add_48_2_groupi_n_1415, csa_tree_add_48_2_groupi_n_1417,
     csa_tree_add_48_2_groupi_n_1418, csa_tree_add_48_2_groupi_n_1419,
     csa_tree_add_48_2_groupi_n_1420, csa_tree_add_48_2_groupi_n_1421,
     csa_tree_add_48_2_groupi_n_1422, csa_tree_add_48_2_groupi_n_1423,
     csa_tree_add_48_2_groupi_n_1424, csa_tree_add_48_2_groupi_n_1425,
     csa_tree_add_48_2_groupi_n_1426, csa_tree_add_48_2_groupi_n_1427,
     csa_tree_add_48_2_groupi_n_1428, csa_tree_add_48_2_groupi_n_1429,
     csa_tree_add_48_2_groupi_n_1430, csa_tree_add_48_2_groupi_n_1431,
     csa_tree_add_48_2_groupi_n_1432, csa_tree_add_48_2_groupi_n_1433,
     csa_tree_add_48_2_groupi_n_1434, csa_tree_add_48_2_groupi_n_1436,
     csa_tree_add_48_2_groupi_n_1437, csa_tree_add_48_2_groupi_n_1438,
     csa_tree_add_48_2_groupi_n_1439, csa_tree_add_48_2_groupi_n_1440,
     csa_tree_add_48_2_groupi_n_1441, csa_tree_add_48_2_groupi_n_1442,
     csa_tree_add_48_2_groupi_n_1443, csa_tree_add_48_2_groupi_n_1444,
     csa_tree_add_48_2_groupi_n_1445, csa_tree_add_48_2_groupi_n_1446,
     csa_tree_add_48_2_groupi_n_1447, csa_tree_add_48_2_groupi_n_1448,
     csa_tree_add_48_2_groupi_n_1449, csa_tree_add_48_2_groupi_n_1450,
     csa_tree_add_48_2_groupi_n_1451, csa_tree_add_48_2_groupi_n_1452,
     csa_tree_add_48_2_groupi_n_1453, csa_tree_add_48_2_groupi_n_1454,
     csa_tree_add_48_2_groupi_n_1455, csa_tree_add_48_2_groupi_n_1456,
     csa_tree_add_48_2_groupi_n_1457, csa_tree_add_48_2_groupi_n_1458,
     csa_tree_add_48_2_groupi_n_1459, csa_tree_add_48_2_groupi_n_1460,
     csa_tree_add_48_2_groupi_n_1461, csa_tree_add_48_2_groupi_n_1462,
     csa_tree_add_48_2_groupi_n_1463, csa_tree_add_48_2_groupi_n_1464,
     csa_tree_add_48_2_groupi_n_1465, csa_tree_add_48_2_groupi_n_1466,
     csa_tree_add_48_2_groupi_n_1467, csa_tree_add_48_2_groupi_n_1468,
     csa_tree_add_48_2_groupi_n_1469, csa_tree_add_48_2_groupi_n_1470,
     csa_tree_add_48_2_groupi_n_1471, csa_tree_add_48_2_groupi_n_1472,
     csa_tree_add_48_2_groupi_n_1473, csa_tree_add_48_2_groupi_n_1474,
     csa_tree_add_48_2_groupi_n_1475, csa_tree_add_48_2_groupi_n_1476,
     csa_tree_add_48_2_groupi_n_1477, csa_tree_add_48_2_groupi_n_1480,
     csa_tree_add_48_2_groupi_n_1481, csa_tree_add_48_2_groupi_n_1482,
     csa_tree_add_48_2_groupi_n_1483, csa_tree_add_48_2_groupi_n_1484,
     csa_tree_add_48_2_groupi_n_1485, csa_tree_add_48_2_groupi_n_1486,
     csa_tree_add_48_2_groupi_n_1487, csa_tree_add_48_2_groupi_n_1488,
     csa_tree_add_48_2_groupi_n_1489, csa_tree_add_48_2_groupi_n_1490,
     csa_tree_add_48_2_groupi_n_1491, csa_tree_add_48_2_groupi_n_1492,
     csa_tree_add_48_2_groupi_n_1493, csa_tree_add_48_2_groupi_n_1494,
     csa_tree_add_48_2_groupi_n_1495, csa_tree_add_48_2_groupi_n_1498,
     csa_tree_add_48_2_groupi_n_1499, csa_tree_add_48_2_groupi_n_1500,
     csa_tree_add_48_2_groupi_n_1501, csa_tree_add_48_2_groupi_n_1502,
     csa_tree_add_48_2_groupi_n_1505, csa_tree_add_48_2_groupi_n_1506,
     csa_tree_add_48_2_groupi_n_1507, csa_tree_add_48_2_groupi_n_1508,
     csa_tree_add_48_2_groupi_n_1510, csa_tree_add_48_2_groupi_n_1511,
     csa_tree_add_48_2_groupi_n_1512, csa_tree_add_48_2_groupi_n_1513,
     csa_tree_add_48_2_groupi_n_1514, csa_tree_add_48_2_groupi_n_1515,
     csa_tree_add_48_2_groupi_n_1516, csa_tree_add_48_2_groupi_n_1517,
     csa_tree_add_48_2_groupi_n_1518, csa_tree_add_48_2_groupi_n_1519,
     csa_tree_add_48_2_groupi_n_1520, csa_tree_add_48_2_groupi_n_1521,
     csa_tree_add_48_2_groupi_n_1522, csa_tree_add_48_2_groupi_n_1523,
     csa_tree_add_48_2_groupi_n_1524, csa_tree_add_48_2_groupi_n_1525,
     csa_tree_add_48_2_groupi_n_1526, csa_tree_add_48_2_groupi_n_1527,
     csa_tree_add_48_2_groupi_n_1528, csa_tree_add_48_2_groupi_n_1529,
     csa_tree_add_48_2_groupi_n_1530, csa_tree_add_48_2_groupi_n_1531,
     csa_tree_add_48_2_groupi_n_1532, csa_tree_add_48_2_groupi_n_1533,
     csa_tree_add_48_2_groupi_n_1534, csa_tree_add_48_2_groupi_n_1535,
     csa_tree_add_48_2_groupi_n_1536, csa_tree_add_48_2_groupi_n_1537,
     csa_tree_add_48_2_groupi_n_1538, csa_tree_add_48_2_groupi_n_1539,
     csa_tree_add_48_2_groupi_n_1540, csa_tree_add_48_2_groupi_n_1541,
     csa_tree_add_48_2_groupi_n_1542, csa_tree_add_48_2_groupi_n_1543,
     csa_tree_add_48_2_groupi_n_1544, csa_tree_add_48_2_groupi_n_1545,
     csa_tree_add_48_2_groupi_n_1546, csa_tree_add_48_2_groupi_n_1547,
     csa_tree_add_48_2_groupi_n_1548, csa_tree_add_48_2_groupi_n_1557,
     csa_tree_add_48_2_groupi_n_1558, csa_tree_add_48_2_groupi_n_1559,
     csa_tree_add_48_2_groupi_n_1560, csa_tree_add_48_2_groupi_n_1561,
     csa_tree_add_48_2_groupi_n_1564, csa_tree_add_48_2_groupi_n_1565,
     csa_tree_add_48_2_groupi_n_1566, csa_tree_add_48_2_groupi_n_1567,
     csa_tree_add_48_2_groupi_n_1570, csa_tree_add_48_2_groupi_n_1571,
     csa_tree_add_48_2_groupi_n_1572, csa_tree_add_48_2_groupi_n_1573,
     csa_tree_add_48_2_groupi_n_1574, csa_tree_add_48_2_groupi_n_1575,
     csa_tree_add_48_2_groupi_n_1576, csa_tree_add_48_2_groupi_n_1577,
     csa_tree_add_48_2_groupi_n_1578, csa_tree_add_48_2_groupi_n_1579,
     csa_tree_add_48_2_groupi_n_1580, csa_tree_add_48_2_groupi_n_1581,
     csa_tree_add_48_2_groupi_n_1582, csa_tree_add_48_2_groupi_n_1583,
     csa_tree_add_48_2_groupi_n_1584, csa_tree_add_48_2_groupi_n_1589,
     csa_tree_add_48_2_groupi_n_1590, csa_tree_add_48_2_groupi_n_1591,
     csa_tree_add_48_2_groupi_n_1592, csa_tree_add_48_2_groupi_n_1593,
     csa_tree_add_48_2_groupi_n_1594, csa_tree_add_48_2_groupi_n_1595,
     csa_tree_add_48_2_groupi_n_1596, csa_tree_add_48_2_groupi_n_1597,
     csa_tree_add_48_2_groupi_n_1598, csa_tree_add_48_2_groupi_n_1600,
     csa_tree_add_48_2_groupi_n_1601, csa_tree_add_48_2_groupi_n_1602,
     csa_tree_add_48_2_groupi_n_1603, csa_tree_add_48_2_groupi_n_1606,
     csa_tree_add_48_2_groupi_n_1607, csa_tree_add_48_2_groupi_n_1608,
     csa_tree_add_48_2_groupi_n_1609, csa_tree_add_48_2_groupi_n_1610,
     csa_tree_add_48_2_groupi_n_1611, csa_tree_add_48_2_groupi_n_1612,
     csa_tree_add_48_2_groupi_n_1613, csa_tree_add_48_2_groupi_n_1614,
     csa_tree_add_48_2_groupi_n_1615, csa_tree_add_48_2_groupi_n_1616,
     csa_tree_add_48_2_groupi_n_1618, csa_tree_add_48_2_groupi_n_1619,
     csa_tree_add_48_2_groupi_n_1620, csa_tree_add_48_2_groupi_n_1621,
     csa_tree_add_48_2_groupi_n_1622, csa_tree_add_48_2_groupi_n_1623,
     csa_tree_add_48_2_groupi_n_1624, csa_tree_add_48_2_groupi_n_1625,
     csa_tree_add_48_2_groupi_n_1626, csa_tree_add_48_2_groupi_n_1627,
     csa_tree_add_48_2_groupi_n_1630, csa_tree_add_48_2_groupi_n_1631,
     csa_tree_add_48_2_groupi_n_1632, csa_tree_add_48_2_groupi_n_1633,
     csa_tree_add_48_2_groupi_n_1634, csa_tree_add_48_2_groupi_n_1635,
     csa_tree_add_48_2_groupi_n_1636, csa_tree_add_48_2_groupi_n_1637,
     csa_tree_add_48_2_groupi_n_1638, csa_tree_add_48_2_groupi_n_1639,
     csa_tree_add_48_2_groupi_n_1640, csa_tree_add_48_2_groupi_n_1646,
     csa_tree_add_48_2_groupi_n_1647, csa_tree_add_48_2_groupi_n_1648,
     csa_tree_add_48_2_groupi_n_1649, csa_tree_add_48_2_groupi_n_1650,
     csa_tree_add_48_2_groupi_n_1651, csa_tree_add_48_2_groupi_n_1652,
     csa_tree_add_48_2_groupi_n_1653, csa_tree_add_48_2_groupi_n_1654,
     csa_tree_add_48_2_groupi_n_1655, csa_tree_add_48_2_groupi_n_1657,
     csa_tree_add_48_2_groupi_n_1659, csa_tree_add_48_2_groupi_n_1660,
     csa_tree_add_48_2_groupi_n_1661, csa_tree_add_48_2_groupi_n_1662,
     csa_tree_add_48_2_groupi_n_1663, csa_tree_add_48_2_groupi_n_1664,
     csa_tree_add_48_2_groupi_n_1665, csa_tree_add_48_2_groupi_n_1666,
     csa_tree_add_48_2_groupi_n_1667, csa_tree_add_48_2_groupi_n_1668,
     csa_tree_add_48_2_groupi_n_1669, csa_tree_add_48_2_groupi_n_1670,
     csa_tree_add_48_2_groupi_n_1671, csa_tree_add_48_2_groupi_n_1672,
     csa_tree_add_48_2_groupi_n_1673, csa_tree_add_48_2_groupi_n_1674,
     csa_tree_add_48_2_groupi_n_1675, csa_tree_add_48_2_groupi_n_1676,
     csa_tree_add_48_2_groupi_n_1677, csa_tree_add_48_2_groupi_n_1678,
     csa_tree_add_48_2_groupi_n_1679, csa_tree_add_48_2_groupi_n_1680,
     csa_tree_add_48_2_groupi_n_1681, csa_tree_add_48_2_groupi_n_1682,
     csa_tree_add_48_2_groupi_n_1683, csa_tree_add_48_2_groupi_n_1684,
     csa_tree_add_48_2_groupi_n_1685, csa_tree_add_48_2_groupi_n_1686,
     csa_tree_add_48_2_groupi_n_1687, csa_tree_add_48_2_groupi_n_1688,
     csa_tree_add_48_2_groupi_n_1689, csa_tree_add_48_2_groupi_n_1690,
     csa_tree_add_48_2_groupi_n_1691, csa_tree_add_48_2_groupi_n_1692,
     csa_tree_add_48_2_groupi_n_1693, csa_tree_add_48_2_groupi_n_1694,
     csa_tree_add_48_2_groupi_n_1695, csa_tree_add_48_2_groupi_n_1696,
     csa_tree_add_48_2_groupi_n_1697, csa_tree_add_48_2_groupi_n_1698,
     csa_tree_add_48_2_groupi_n_1699, csa_tree_add_48_2_groupi_n_1700,
     csa_tree_add_48_2_groupi_n_1701, csa_tree_add_48_2_groupi_n_1702,
     csa_tree_add_48_2_groupi_n_1703, csa_tree_add_48_2_groupi_n_1704,
     csa_tree_add_48_2_groupi_n_1705, csa_tree_add_48_2_groupi_n_1706,
     csa_tree_add_48_2_groupi_n_1707, csa_tree_add_48_2_groupi_n_1708,
     csa_tree_add_48_2_groupi_n_1709, csa_tree_add_48_2_groupi_n_1710,
     csa_tree_add_48_2_groupi_n_1711, csa_tree_add_48_2_groupi_n_1712,
     csa_tree_add_48_2_groupi_n_1713, csa_tree_add_48_2_groupi_n_1714,
     csa_tree_add_48_2_groupi_n_1715, csa_tree_add_48_2_groupi_n_1716,
     csa_tree_add_48_2_groupi_n_1718, csa_tree_add_48_2_groupi_n_1719,
     csa_tree_add_48_2_groupi_n_1720, csa_tree_add_48_2_groupi_n_1721,
     csa_tree_add_48_2_groupi_n_1722, csa_tree_add_48_2_groupi_n_1723,
     csa_tree_add_48_2_groupi_n_1724, csa_tree_add_48_2_groupi_n_1725,
     csa_tree_add_48_2_groupi_n_1726, csa_tree_add_48_2_groupi_n_1727,
     csa_tree_add_48_2_groupi_n_1728, csa_tree_add_48_2_groupi_n_1729,
     csa_tree_add_48_2_groupi_n_1731, csa_tree_add_48_2_groupi_n_1732,
     csa_tree_add_48_2_groupi_n_1733, csa_tree_add_48_2_groupi_n_1734,
     csa_tree_add_48_2_groupi_n_1736, csa_tree_add_48_2_groupi_n_1737,
     csa_tree_add_48_2_groupi_n_1738, csa_tree_add_48_2_groupi_n_1740,
     csa_tree_add_48_2_groupi_n_1741, csa_tree_add_48_2_groupi_n_1742,
     csa_tree_add_48_2_groupi_n_1744, csa_tree_add_48_2_groupi_n_1745,
     csa_tree_add_48_2_groupi_n_1746, csa_tree_add_48_2_groupi_n_1747,
     csa_tree_add_48_2_groupi_n_1748, csa_tree_add_48_2_groupi_n_1750,
     csa_tree_add_48_2_groupi_n_1751, csa_tree_add_48_2_groupi_n_1752,
     csa_tree_add_48_2_groupi_n_1754, csa_tree_add_48_2_groupi_n_1755,
     csa_tree_add_48_2_groupi_n_1756, csa_tree_add_48_2_groupi_n_1758,
     csa_tree_add_48_2_groupi_n_1759, csa_tree_add_48_2_groupi_n_1760,
     csa_tree_add_48_2_groupi_n_1762, csa_tree_add_48_2_groupi_n_1763,
     csa_tree_add_48_2_groupi_n_1764, csa_tree_add_48_2_groupi_n_1766,
     csa_tree_add_48_2_groupi_n_1767, csa_tree_add_48_2_groupi_n_1769,
     csa_tree_add_48_2_groupi_n_1770, csa_tree_add_48_2_groupi_n_1771,
     csa_tree_add_48_2_groupi_n_1773, csa_tree_add_48_2_groupi_n_1774,
     csa_tree_add_48_2_groupi_n_1775, csa_tree_add_48_2_groupi_n_1777,
     csa_tree_add_48_2_groupi_n_1779, n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7,
     n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20,
     n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31, n_32,
     n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_41, n_42, n_43, n_44,
     n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55, n_56,
     n_57, n_58, n_59, n_60, clk, n_164, n_165, n_166, n_167, n_168, n_169,
     n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180,
     n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188, n_189;
 reg out1_7_L0_reg_N30;
 always @(posedge clk)
         out1_7_L0_reg_N30 <= n_19;
 assign {out1[24]} = out1_7_L0_reg_N30;
 reg out1_8_L0_reg_N30;
 always @(posedge clk)
         out1_8_L0_reg_N30 <= n_23;
 assign {out1[23]} = out1_8_L0_reg_N30;
 reg out1_9_L0_reg_N30;
 always @(posedge clk)
         out1_9_L0_reg_N30 <= n_40;
 assign {out1[22]} = out1_9_L0_reg_N30;
 reg out1_10_L0_reg_N30;
 always @(posedge clk)
         out1_10_L0_reg_N30 <= n_44;
 assign {out1[21]} = out1_10_L0_reg_N30;
 reg out1_11_L0_reg_N30;
 always @(posedge clk)
         out1_11_L0_reg_N30 <= n_47;
 assign {out1[20]} = out1_11_L0_reg_N30;
 reg out1_12_L0_reg_N30;
 always @(posedge clk)
         out1_12_L0_reg_N30 <= n_54;
 assign {out1[19]} = out1_12_L0_reg_N30;
 reg out1_13_L0_reg_N30;
 always @(posedge clk)
         out1_13_L0_reg_N30 <= n_49;
 assign {out1[18]} = out1_13_L0_reg_N30;
 reg out1_14_L0_reg_N30;
 always @(posedge clk)
         out1_14_L0_reg_N30 <= n_48;
 assign {out1[17]} = out1_14_L0_reg_N30;
 reg out1_15_L0_reg_N30;
 always @(posedge clk)
         out1_15_L0_reg_N30 <= n_43;
 assign {out1[16]} = out1_15_L0_reg_N30;
 reg out1_16_L0_reg_N30;
 always @(posedge clk)
         out1_16_L0_reg_N30 <= n_53;
 assign {out1[15]} = out1_16_L0_reg_N30;
 reg out1_17_L0_reg_N30;
 always @(posedge clk)
         out1_17_L0_reg_N30 <= n_52;
 assign {out1[14]} = out1_17_L0_reg_N30;
 reg out1_18_L0_reg_N30;
 always @(posedge clk)
         out1_18_L0_reg_N30 <= n_46;
 assign {out1[13]} = out1_18_L0_reg_N30;
 reg out1_19_L0_reg_N30;
 always @(posedge clk)
         if (csa_tree_add_48_2_groupi_n_1744)
         out1_19_L0_reg_N30 <= n_56;
     else
         out1_19_L0_reg_N30 <= csa_tree_add_48_2_groupi_n_107;
 assign {out1[12]} = out1_19_L0_reg_N30;
 reg out1_20_L0_reg_N30;
 always @(posedge clk)
         out1_20_L0_reg_N30 <= n_42;
 assign {out1[11]} = out1_20_L0_reg_N30;
 reg out1_21_L0_reg_N30;
 always @(posedge clk)
         out1_21_L0_reg_N30 <= n_55;
 assign {out1[10]} = out1_21_L0_reg_N30;
 reg out1_22_L0_reg_N30;
 always @(posedge clk)
         out1_22_L0_reg_N30 <= n_50;
 assign {out1[9]} = out1_22_L0_reg_N30;
 reg out1_23_L0_reg_N30;
 always @(posedge clk)
         out1_23_L0_reg_N30 <= n_51;
 assign {out1[8]} = out1_23_L0_reg_N30;
 reg out1_24_L0_reg_N30;
 always @(posedge clk)
         out1_24_L0_reg_N30 <= n_45;
 assign {out1[7]} = out1_24_L0_reg_N30;
 reg out1_25_L0_reg_N30;
 always @(posedge clk)
         if (csa_tree_add_48_2_groupi_n_1637)
         out1_25_L0_reg_N30 <= n_58;
     else
         out1_25_L0_reg_N30 <= csa_tree_add_48_2_groupi_n_1657;
 assign {out1[6]} = out1_25_L0_reg_N30;
 reg out1_26_L0_reg_N30;
 always @(posedge clk)
         if (csa_tree_add_48_2_groupi_n_1619)
         out1_26_L0_reg_N30 <= n_57;
     else
         out1_26_L0_reg_N30 <= csa_tree_add_48_2_groupi_n_1625;
 assign {out1[5]} = out1_26_L0_reg_N30;
 reg out1_27_L0_reg_N30;
 always @(posedge clk)
         if (csa_tree_add_48_2_groupi_n_1578)
         out1_27_L0_reg_N30 <= n_59;
     else
         out1_27_L0_reg_N30 <= csa_tree_add_48_2_groupi_n_1543;
 assign {out1[4]} = out1_27_L0_reg_N30;
 reg out1_28_L0_reg_N30;
 always @(posedge clk)
         if (csa_tree_add_48_2_groupi_n_1495)
         out1_28_L0_reg_N30 <= n_60;
     else
         out1_28_L0_reg_N30 <= csa_tree_add_48_2_groupi_n_1499;
 assign {out1[3]} = out1_28_L0_reg_N30;
 reg out1_29_L0_reg_N30;
 always @(posedge clk)
         out1_29_L0_reg_N30 <= n_21;
 assign {out1[2]} = out1_29_L0_reg_N30;
 reg out1_30_L0_reg_N30;
 always @(posedge clk)
         out1_30_L0_reg_N30 <= n_22;
 assign {out1[1]} = out1_30_L0_reg_N30;
 reg out1_31_L0_reg_N30;
 always @(posedge clk)
         out1_31_L0_reg_N30 <= n_34;
 assign {out1[0]} = out1_31_L0_reg_N30;
 reg retime_s1_1_reg_reg_N30;
 always @(posedge clk)
         retime_s1_1_reg_reg_N30 <= n_18;
 assign n_0 = retime_s1_1_reg_reg_N30;
 reg retime_s1_2_reg_reg_N30;
 always @(posedge clk)
         retime_s1_2_reg_reg_N30 <= n_17;
 assign {out1[25]} = retime_s1_2_reg_reg_N30;
 reg retime_s1_3_reg_reg_N30;
 always @(posedge clk)
         retime_s1_3_reg_reg_N30 <= n_29;
 assign n_1 = retime_s1_3_reg_reg_N30;
 reg retime_s1_4_reg_reg_N30;
 always @(posedge clk)
         retime_s1_4_reg_reg_N30 <= n_37;
 assign n_2 = retime_s1_4_reg_reg_N30;
 reg retime_s1_5_reg_reg_N30;
 always @(posedge clk)
         retime_s1_5_reg_reg_N30 <= n_36;
 assign n_3 = retime_s1_5_reg_reg_N30;
 reg retime_s1_6_reg_reg_N30;
 always @(posedge clk)
         retime_s1_6_reg_reg_N30 <= n_33;
 assign n_4 = retime_s1_6_reg_reg_N30;
 reg retime_s1_7_reg_reg_N30;
 always @(posedge clk)
         retime_s1_7_reg_reg_N30 <= n_32;
 assign n_5 = retime_s1_7_reg_reg_N30;
 reg retime_s1_8_reg_reg_N30;
 always @(posedge clk)
         retime_s1_8_reg_reg_N30 <= n_39;
 assign n_6 = retime_s1_8_reg_reg_N30;
 reg retime_s1_9_reg_reg_N30;
 always @(posedge clk)
         retime_s1_9_reg_reg_N30 <= n_38;
 assign n_7 = retime_s1_9_reg_reg_N30;
 reg retime_s1_10_reg_reg_N30;
 always @(posedge clk)
         retime_s1_10_reg_reg_N30 <= n_27;
 assign n_8 = retime_s1_10_reg_reg_N30;
 reg retime_s1_11_reg_reg_N30;
 always @(posedge clk)
         retime_s1_11_reg_reg_N30 <= n_26;
 assign n_9 = retime_s1_11_reg_reg_N30;
 reg retime_s1_12_reg_reg_N30;
 always @(posedge clk)
         retime_s1_12_reg_reg_N30 <= n_30;
 assign n_10 = retime_s1_12_reg_reg_N30;
 reg retime_s1_13_reg_reg_N30;
 always @(posedge clk)
         retime_s1_13_reg_reg_N30 <= n_25;
 assign n_11 = retime_s1_13_reg_reg_N30;
 assign csa_tree_add_48_2_groupi_n_115 = ({in2[7]} & {in1[0]});
 assign csa_tree_add_48_2_groupi_n_1779 = ~(csa_tree_add_48_2_groupi_n_1580 & (csa_tree_add_48_2_groupi_n_1777
    | csa_tree_add_48_2_groupi_n_1612));
 assign csa_tree_add_48_2_groupi_n_1777 = ~(csa_tree_add_48_2_groupi_n_1775 | csa_tree_add_48_2_groupi_n_1597);
 assign csa_tree_add_48_2_groupi_n_1775 = ~(csa_tree_add_48_2_groupi_n_1773 | csa_tree_add_48_2_groupi_n_1603);
 assign csa_tree_add_48_2_groupi_n_1774 = ~csa_tree_add_48_2_groupi_n_1773;
 assign csa_tree_add_48_2_groupi_n_1773 = ~(csa_tree_add_48_2_groupi_n_1771 | csa_tree_add_48_2_groupi_n_1659);
 assign csa_tree_add_48_2_groupi_n_1771 = ~(csa_tree_add_48_2_groupi_n_1769 | csa_tree_add_48_2_groupi_n_1664);
 assign csa_tree_add_48_2_groupi_n_1770 = ~csa_tree_add_48_2_groupi_n_1769;
 assign csa_tree_add_48_2_groupi_n_1769 = ~(csa_tree_add_48_2_groupi_n_1767 | csa_tree_add_48_2_groupi_n_1685);
 assign csa_tree_add_48_2_groupi_n_1767 = ~(csa_tree_add_48_2_groupi_n_1688 | ~(csa_tree_add_48_2_groupi_n_1764
    | csa_tree_add_48_2_groupi_n_1684));
 assign csa_tree_add_48_2_groupi_n_1766 = (csa_tree_add_48_2_groupi_n_1764 | csa_tree_add_48_2_groupi_n_1684);
 assign csa_tree_add_48_2_groupi_n_1764 = ~(csa_tree_add_48_2_groupi_n_1762 | csa_tree_add_48_2_groupi_n_1687);
 assign csa_tree_add_48_2_groupi_n_1763 = ~csa_tree_add_48_2_groupi_n_1762;
 assign csa_tree_add_48_2_groupi_n_1762 = ~(csa_tree_add_48_2_groupi_n_1760 | ~csa_tree_add_48_2_groupi_n_1699);
 assign csa_tree_add_48_2_groupi_n_1760 = ~(csa_tree_add_48_2_groupi_n_1758 | csa_tree_add_48_2_groupi_n_1701);
 assign csa_tree_add_48_2_groupi_n_1759 = ~csa_tree_add_48_2_groupi_n_1758;
 assign csa_tree_add_48_2_groupi_n_1758 = ~(csa_tree_add_48_2_groupi_n_1756 | csa_tree_add_48_2_groupi_n_1700);
 assign csa_tree_add_48_2_groupi_n_1756 = ~(csa_tree_add_48_2_groupi_n_1754 | csa_tree_add_48_2_groupi_n_1703);
 assign csa_tree_add_48_2_groupi_n_1755 = ~csa_tree_add_48_2_groupi_n_1754;
 assign csa_tree_add_48_2_groupi_n_1754 = ~(csa_tree_add_48_2_groupi_n_1752 | csa_tree_add_48_2_groupi_n_1713);
 assign csa_tree_add_48_2_groupi_n_1752 = ~(csa_tree_add_48_2_groupi_n_1750 | ~csa_tree_add_48_2_groupi_n_1715);
 assign csa_tree_add_48_2_groupi_n_1751 = ~csa_tree_add_48_2_groupi_n_1750;
 assign csa_tree_add_48_2_groupi_n_1750 = ~(csa_tree_add_48_2_groupi_n_1748 | csa_tree_add_48_2_groupi_n_1727);
 assign csa_tree_add_48_2_groupi_n_1748 = ~(csa_tree_add_48_2_groupi_n_1746 | ~csa_tree_add_48_2_groupi_n_1728);
 assign csa_tree_add_48_2_groupi_n_1747 = ~csa_tree_add_48_2_groupi_n_1746;
 assign csa_tree_add_48_2_groupi_n_1746 = ~(csa_tree_add_48_2_groupi_n_1745 | csa_tree_add_48_2_groupi_n_1726);
 assign csa_tree_add_48_2_groupi_n_1745 = ~(csa_tree_add_48_2_groupi_n_1744 | ~csa_tree_add_48_2_groupi_n_1729);
 assign csa_tree_add_48_2_groupi_n_1744 = ~(csa_tree_add_48_2_groupi_n_1742 | ~csa_tree_add_48_2_groupi_n_1716);
 assign csa_tree_add_48_2_groupi_n_1742 = ~(csa_tree_add_48_2_groupi_n_1740 | ~csa_tree_add_48_2_groupi_n_1714);
 assign csa_tree_add_48_2_groupi_n_1741 = ~csa_tree_add_48_2_groupi_n_1740;
 assign csa_tree_add_48_2_groupi_n_1740 = ~(csa_tree_add_48_2_groupi_n_1738 | ~csa_tree_add_48_2_groupi_n_1698);
 assign csa_tree_add_48_2_groupi_n_1738 = ~(csa_tree_add_48_2_groupi_n_1736 | ~csa_tree_add_48_2_groupi_n_1702);
 assign csa_tree_add_48_2_groupi_n_1737 = ~csa_tree_add_48_2_groupi_n_1736;
 assign csa_tree_add_48_2_groupi_n_1736 = ~(csa_tree_add_48_2_groupi_n_1734 | csa_tree_add_48_2_groupi_n_106);
 assign csa_tree_add_48_2_groupi_n_1734 = ~(csa_tree_add_48_2_groupi_n_1731 | csa_tree_add_48_2_groupi_n_1686);
 assign csa_tree_add_48_2_groupi_n_1733 = ~csa_tree_add_48_2_groupi_n_1731;
 assign csa_tree_add_48_2_groupi_n_1732 = ~(csa_tree_add_48_2_groupi_n_1707 ^ csa_tree_add_48_2_groupi_n_1720);
 assign csa_tree_add_48_2_groupi_n_1731 = ~(csa_tree_add_48_2_groupi_n_1725 | ~csa_tree_add_48_2_groupi_n_1668);
 assign csa_tree_add_48_2_groupi_n_1729 = ~(csa_tree_add_48_2_groupi_n_1718 & ~csa_tree_add_48_2_groupi_n_1673);
 assign csa_tree_add_48_2_groupi_n_1728 = ~(csa_tree_add_48_2_groupi_n_1708 & csa_tree_add_48_2_groupi_n_1723);
 assign csa_tree_add_48_2_groupi_n_1727 = ~(csa_tree_add_48_2_groupi_n_1708 | csa_tree_add_48_2_groupi_n_1723);
 assign csa_tree_add_48_2_groupi_n_1726 = ~(csa_tree_add_48_2_groupi_n_1718 | ~csa_tree_add_48_2_groupi_n_1673);
 assign csa_tree_add_48_2_groupi_n_1725 = ~(csa_tree_add_48_2_groupi_n_1719 | ~csa_tree_add_48_2_groupi_n_1669);
 assign csa_tree_add_48_2_groupi_n_1724 = ~csa_tree_add_48_2_groupi_n_1719;
 assign csa_tree_add_48_2_groupi_n_1723 = ~csa_tree_add_48_2_groupi_n_1720;
 assign csa_tree_add_48_2_groupi_n_1722 = ~(csa_tree_add_48_2_groupi_n_1690 ^ csa_tree_add_48_2_groupi_n_1706);
 assign csa_tree_add_48_2_groupi_n_1721 = ~(csa_tree_add_48_2_groupi_n_1691 ^ csa_tree_add_48_2_groupi_n_1705);
 assign csa_tree_add_48_2_groupi_n_1720 = ~(csa_tree_add_48_2_groupi_n_1675 & (csa_tree_add_48_2_groupi_n_1676
    | csa_tree_add_48_2_groupi_n_1652));
 assign csa_tree_add_48_2_groupi_n_1719 = ~(csa_tree_add_48_2_groupi_n_1712 | ~csa_tree_add_48_2_groupi_n_1638);
 assign csa_tree_add_48_2_groupi_n_1718 = ~((csa_tree_add_48_2_groupi_n_1652 & ~csa_tree_add_48_2_groupi_n_99)
    | (csa_tree_add_48_2_groupi_n_1651 & csa_tree_add_48_2_groupi_n_99));
 assign csa_tree_add_48_2_groupi_n_1716 = ~(csa_tree_add_48_2_groupi_n_1705 & csa_tree_add_48_2_groupi_n_1691);
 assign csa_tree_add_48_2_groupi_n_1715 = (csa_tree_add_48_2_groupi_n_1690 | csa_tree_add_48_2_groupi_n_1706);
 assign csa_tree_add_48_2_groupi_n_1714 = ~(csa_tree_add_48_2_groupi_n_103 & csa_tree_add_48_2_groupi_n_1672);
 assign csa_tree_add_48_2_groupi_n_1713 = (csa_tree_add_48_2_groupi_n_1690 & csa_tree_add_48_2_groupi_n_1706);
 assign csa_tree_add_48_2_groupi_n_1712 = ~(csa_tree_add_48_2_groupi_n_1683 | csa_tree_add_48_2_groupi_n_1646);
 assign csa_tree_add_48_2_groupi_n_1711 = ~(csa_tree_add_48_2_groupi_n_1680 ^ csa_tree_add_48_2_groupi_n_1693);
 assign csa_tree_add_48_2_groupi_n_1710 = ~(csa_tree_add_48_2_groupi_n_1694 ^ csa_tree_add_48_2_groupi_n_1689);
 assign csa_tree_add_48_2_groupi_n_1709 = ~(csa_tree_add_48_2_groupi_n_1692 ^ csa_tree_add_48_2_groupi_n_1677);
 assign csa_tree_add_48_2_groupi_n_1708 = ~csa_tree_add_48_2_groupi_n_1707;
 assign csa_tree_add_48_2_groupi_n_1705 = ~csa_tree_add_48_2_groupi_n_103;
 assign csa_tree_add_48_2_groupi_n_1704 = ~csa_tree_add_48_2_groupi_n_1683;
 assign csa_tree_add_48_2_groupi_n_1706 = ((csa_tree_add_48_2_groupi_n_1654 & csa_tree_add_48_2_groupi_n_1589)
    | ((csa_tree_add_48_2_groupi_n_1589 & csa_tree_add_48_2_groupi_n_1632) | (csa_tree_add_48_2_groupi_n_1632
    & csa_tree_add_48_2_groupi_n_1654)));
 assign csa_tree_add_48_2_groupi_n_1707 = (csa_tree_add_48_2_groupi_n_1589 ^ (csa_tree_add_48_2_groupi_n_1632
    ^ csa_tree_add_48_2_groupi_n_1654));
 assign csa_tree_add_48_2_groupi_n_1703 = ~(csa_tree_add_48_2_groupi_n_1694 | csa_tree_add_48_2_groupi_n_1689);
 assign csa_tree_add_48_2_groupi_n_1702 = ~(csa_tree_add_48_2_groupi_n_104 & ~csa_tree_add_48_2_groupi_n_1677);
 assign csa_tree_add_48_2_groupi_n_1701 = ~(csa_tree_add_48_2_groupi_n_1693 | csa_tree_add_48_2_groupi_n_1680);
 assign csa_tree_add_48_2_groupi_n_1700 = (csa_tree_add_48_2_groupi_n_1694 & csa_tree_add_48_2_groupi_n_1689);
 assign csa_tree_add_48_2_groupi_n_1699 = ~(csa_tree_add_48_2_groupi_n_1693 & csa_tree_add_48_2_groupi_n_1680);
 assign csa_tree_add_48_2_groupi_n_1698 = ~(csa_tree_add_48_2_groupi_n_1677 & csa_tree_add_48_2_groupi_n_1692);
 assign csa_tree_add_48_2_groupi_n_1697 = ~(csa_tree_add_48_2_groupi_n_1681 ^ csa_tree_add_48_2_groupi_n_1648);
 assign csa_tree_add_48_2_groupi_n_1696 = ~(csa_tree_add_48_2_groupi_n_1679 ^ csa_tree_add_48_2_groupi_n_1682);
 assign csa_tree_add_48_2_groupi_n_1695 = ~(csa_tree_add_48_2_groupi_n_1678 ^ csa_tree_add_48_2_groupi_n_1665);
 assign csa_tree_add_48_2_groupi_n_1692 = ~csa_tree_add_48_2_groupi_n_104;
 assign csa_tree_add_48_2_groupi_n_1691 = ~csa_tree_add_48_2_groupi_n_1672;
 assign csa_tree_add_48_2_groupi_n_1693 = ((csa_tree_add_48_2_groupi_n_1621 & csa_tree_add_48_2_groupi_n_1558)
    | ((csa_tree_add_48_2_groupi_n_1558 & csa_tree_add_48_2_groupi_n_1624) | (csa_tree_add_48_2_groupi_n_1624
    & csa_tree_add_48_2_groupi_n_1621)));
 assign csa_tree_add_48_2_groupi_n_1694 = (csa_tree_add_48_2_groupi_n_1558 ^ (csa_tree_add_48_2_groupi_n_1624
    ^ csa_tree_add_48_2_groupi_n_1621));
 assign csa_tree_add_48_2_groupi_n_1689 = ((csa_tree_add_48_2_groupi_n_1631 & csa_tree_add_48_2_groupi_n_1582)
    | ((csa_tree_add_48_2_groupi_n_1582 & csa_tree_add_48_2_groupi_n_1622) | (csa_tree_add_48_2_groupi_n_1622
    & csa_tree_add_48_2_groupi_n_1631)));
 assign csa_tree_add_48_2_groupi_n_1690 = (csa_tree_add_48_2_groupi_n_1582 ^ (csa_tree_add_48_2_groupi_n_1622
    ^ csa_tree_add_48_2_groupi_n_1631));
 assign csa_tree_add_48_2_groupi_n_1688 = ~(csa_tree_add_48_2_groupi_n_1681 | csa_tree_add_48_2_groupi_n_1648);
 assign csa_tree_add_48_2_groupi_n_1687 = ~(csa_tree_add_48_2_groupi_n_1679 | csa_tree_add_48_2_groupi_n_1682);
 assign csa_tree_add_48_2_groupi_n_1686 = ~(csa_tree_add_48_2_groupi_n_1678 | ~csa_tree_add_48_2_groupi_n_1640);
 assign csa_tree_add_48_2_groupi_n_1685 = (csa_tree_add_48_2_groupi_n_1681 & csa_tree_add_48_2_groupi_n_1648);
 assign csa_tree_add_48_2_groupi_n_1684 = (csa_tree_add_48_2_groupi_n_1679 & csa_tree_add_48_2_groupi_n_1682);
 assign csa_tree_add_48_2_groupi_n_1683 = ~(csa_tree_add_48_2_groupi_n_1674 | ~csa_tree_add_48_2_groupi_n_1627);
 assign csa_tree_add_48_2_groupi_n_1681 = ((csa_tree_add_48_2_groupi_n_1607 & csa_tree_add_48_2_groupi_n_1428)
    | ((csa_tree_add_48_2_groupi_n_1428 & csa_tree_add_48_2_groupi_n_1610) | (csa_tree_add_48_2_groupi_n_1610
    & csa_tree_add_48_2_groupi_n_1607)));
 assign csa_tree_add_48_2_groupi_n_1682 = (csa_tree_add_48_2_groupi_n_1428 ^ (csa_tree_add_48_2_groupi_n_1610
    ^ csa_tree_add_48_2_groupi_n_1607));
 assign csa_tree_add_48_2_groupi_n_1679 = ((csa_tree_add_48_2_groupi_n_1623 & csa_tree_add_48_2_groupi_n_1571)
    | ((csa_tree_add_48_2_groupi_n_1571 & csa_tree_add_48_2_groupi_n_1608) | (csa_tree_add_48_2_groupi_n_1608
    & csa_tree_add_48_2_groupi_n_1623)));
 assign csa_tree_add_48_2_groupi_n_1680 = (csa_tree_add_48_2_groupi_n_1571 ^ (csa_tree_add_48_2_groupi_n_1608
    ^ csa_tree_add_48_2_groupi_n_1623));
 assign csa_tree_add_48_2_groupi_n_1677 = ((csa_tree_add_48_2_groupi_n_1577 & csa_tree_add_48_2_groupi_n_1616)
    | ((csa_tree_add_48_2_groupi_n_1616 & csa_tree_add_48_2_groupi_n_92) | (csa_tree_add_48_2_groupi_n_92
    & csa_tree_add_48_2_groupi_n_1577)));
 assign csa_tree_add_48_2_groupi_n_1678 = (csa_tree_add_48_2_groupi_n_1616 ^ (csa_tree_add_48_2_groupi_n_92
    ^ csa_tree_add_48_2_groupi_n_1577));
 assign csa_tree_add_48_2_groupi_n_1676 = ~(csa_tree_add_48_2_groupi_n_1670 | csa_tree_add_48_2_groupi_n_1591);
 assign csa_tree_add_48_2_groupi_n_1675 = ~(csa_tree_add_48_2_groupi_n_1670 & csa_tree_add_48_2_groupi_n_1591);
 assign csa_tree_add_48_2_groupi_n_1674 = ~(csa_tree_add_48_2_groupi_n_1657 | csa_tree_add_48_2_groupi_n_1630);
 assign csa_tree_add_48_2_groupi_n_1671 = ~(csa_tree_add_48_2_groupi_n_1666 ^ csa_tree_add_48_2_groupi_n_1618);
 assign csa_tree_add_48_2_groupi_n_1673 = ~(csa_tree_add_48_2_groupi_n_1663 & (csa_tree_add_48_2_groupi_n_1662
    | csa_tree_add_48_2_groupi_n_1649));
 assign csa_tree_add_48_2_groupi_n_1672 = ~(csa_tree_add_48_2_groupi_n_1660 | (csa_tree_add_48_2_groupi_n_1661
    & csa_tree_add_48_2_groupi_n_1636));
 assign csa_tree_add_48_2_groupi_n_1670 = ~n_165;
 assign csa_tree_add_48_2_groupi_n_1669 = ~(n_166 & ~csa_tree_add_48_2_groupi_n_1618);
 assign csa_tree_add_48_2_groupi_n_1668 = ~(csa_tree_add_48_2_groupi_n_1666 & csa_tree_add_48_2_groupi_n_1618);
 assign csa_tree_add_48_2_groupi_n_1667 = ~(csa_tree_add_48_2_groupi_n_1596 ^ csa_tree_add_48_2_groupi_n_1647);
 assign csa_tree_add_48_2_groupi_n_1666 = ~n_166;
 assign csa_tree_add_48_2_groupi_n_1665 = ~csa_tree_add_48_2_groupi_n_1640;
 assign csa_tree_add_48_2_groupi_n_1664 = ~(csa_tree_add_48_2_groupi_n_1596 | csa_tree_add_48_2_groupi_n_1647);
 assign csa_tree_add_48_2_groupi_n_1663 = ~(csa_tree_add_48_2_groupi_n_1653 & csa_tree_add_48_2_groupi_n_1635);
 assign csa_tree_add_48_2_groupi_n_1662 = ~(csa_tree_add_48_2_groupi_n_1653 | csa_tree_add_48_2_groupi_n_1635);
 assign csa_tree_add_48_2_groupi_n_1661 = ~(csa_tree_add_48_2_groupi_n_1650 & ~csa_tree_add_48_2_groupi_n_1615);
 assign csa_tree_add_48_2_groupi_n_1660 = ~(csa_tree_add_48_2_groupi_n_1650 | ~csa_tree_add_48_2_groupi_n_1615);
 assign csa_tree_add_48_2_groupi_n_1659 = (csa_tree_add_48_2_groupi_n_1596 & csa_tree_add_48_2_groupi_n_1647);
 assign csa_tree_add_48_2_groupi_n_1655 = ~(n_167 ^ csa_tree_add_48_2_groupi_n_1600);
 assign csa_tree_add_48_2_groupi_n_1654 = ~(csa_tree_add_48_2_groupi_n_1542 & (csa_tree_add_48_2_groupi_n_1634
    | csa_tree_add_48_2_groupi_n_1545));
 assign csa_tree_add_48_2_groupi_n_1657 = ~(csa_tree_add_48_2_groupi_n_1639 | csa_tree_add_48_2_groupi_n_100);
 assign csa_tree_add_48_2_groupi_n_1652 = ~csa_tree_add_48_2_groupi_n_1651;
 assign csa_tree_add_48_2_groupi_n_1651 = ((csa_tree_add_48_2_groupi_n_1611 & csa_tree_add_48_2_groupi_n_1492)
    | ((csa_tree_add_48_2_groupi_n_1492 & csa_tree_add_48_2_groupi_n_1530) | (csa_tree_add_48_2_groupi_n_1530
    & csa_tree_add_48_2_groupi_n_1611)));
 assign csa_tree_add_48_2_groupi_n_1653 = (csa_tree_add_48_2_groupi_n_1492 ^ (csa_tree_add_48_2_groupi_n_1530
    ^ csa_tree_add_48_2_groupi_n_1611));
 assign csa_tree_add_48_2_groupi_n_1649 = ((csa_tree_add_48_2_groupi_n_1541 & csa_tree_add_48_2_groupi_n_1521)
    | ((csa_tree_add_48_2_groupi_n_1521 & csa_tree_add_48_2_groupi_n_84) | (csa_tree_add_48_2_groupi_n_84
    & csa_tree_add_48_2_groupi_n_1541)));
 assign csa_tree_add_48_2_groupi_n_1650 = (csa_tree_add_48_2_groupi_n_1521 ^ (csa_tree_add_48_2_groupi_n_84
    ^ csa_tree_add_48_2_groupi_n_1541));
 assign csa_tree_add_48_2_groupi_n_1647 = ((csa_tree_add_48_2_groupi_n_1609 & csa_tree_add_48_2_groupi_n_1427)
    | ((csa_tree_add_48_2_groupi_n_1427 & csa_tree_add_48_2_groupi_n_1512) | (csa_tree_add_48_2_groupi_n_1512
    & csa_tree_add_48_2_groupi_n_1609)));
 assign csa_tree_add_48_2_groupi_n_1648 = (csa_tree_add_48_2_groupi_n_1427 ^ (csa_tree_add_48_2_groupi_n_1512
    ^ csa_tree_add_48_2_groupi_n_1609));
 assign csa_tree_add_48_2_groupi_n_1646 = ~(n_167 | csa_tree_add_48_2_groupi_n_1600);
 assign csa_tree_add_48_2_groupi_n_1639 = ~(csa_tree_add_48_2_groupi_n_1625 | csa_tree_add_48_2_groupi_n_1602);
 assign csa_tree_add_48_2_groupi_n_1638 = ~(n_167 & csa_tree_add_48_2_groupi_n_1600);
 assign csa_tree_add_48_2_groupi_n_1637 = ~(n_168 ^ csa_tree_add_48_2_groupi_n_1593);
 assign csa_tree_add_48_2_groupi_n_1640 = ~(csa_tree_add_48_2_groupi_n_1626 | csa_tree_add_48_2_groupi_n_1606);
 assign csa_tree_add_48_2_groupi_n_1636 = ~csa_tree_add_48_2_groupi_n_1584;
 assign csa_tree_add_48_2_groupi_n_1634 = ~csa_tree_add_48_2_groupi_n_1633;
 assign csa_tree_add_48_2_groupi_n_1631 = ((csa_tree_add_48_2_groupi_n_1473 & csa_tree_add_48_2_groupi_n_1583)
    | ((csa_tree_add_48_2_groupi_n_1583 & csa_tree_add_48_2_groupi_n_1514) | (csa_tree_add_48_2_groupi_n_1514
    & csa_tree_add_48_2_groupi_n_1473)));
 assign csa_tree_add_48_2_groupi_n_1632 = (csa_tree_add_48_2_groupi_n_1583 ^ (csa_tree_add_48_2_groupi_n_1514
    ^ csa_tree_add_48_2_groupi_n_1473));
 assign csa_tree_add_48_2_groupi_n_1633 = ((csa_tree_add_48_2_groupi_n_1382 & csa_tree_add_48_2_groupi_n_1510)
    | ((csa_tree_add_48_2_groupi_n_1510 & csa_tree_add_48_2_groupi_n_1493) | (csa_tree_add_48_2_groupi_n_1493
    & csa_tree_add_48_2_groupi_n_1382)));
 assign csa_tree_add_48_2_groupi_n_1635 = (csa_tree_add_48_2_groupi_n_1510 ^ (csa_tree_add_48_2_groupi_n_1493
    ^ csa_tree_add_48_2_groupi_n_1382));
 assign csa_tree_add_48_2_groupi_n_1630 = ~(n_168 | csa_tree_add_48_2_groupi_n_1593);
 assign csa_tree_add_48_2_groupi_n_1627 = ~(n_168 & csa_tree_add_48_2_groupi_n_1593);
 assign csa_tree_add_48_2_groupi_n_1626 = ~(csa_tree_add_48_2_groupi_n_1601 | csa_tree_add_48_2_groupi_n_1581);
 assign csa_tree_add_48_2_groupi_n_1623 = ((csa_tree_add_48_2_groupi_n_1488 & csa_tree_add_48_2_groupi_n_1567)
    | ((csa_tree_add_48_2_groupi_n_1567 & csa_tree_add_48_2_groupi_n_1445) | (csa_tree_add_48_2_groupi_n_1445
    & csa_tree_add_48_2_groupi_n_1488)));
 assign csa_tree_add_48_2_groupi_n_1624 = (csa_tree_add_48_2_groupi_n_1567 ^ (csa_tree_add_48_2_groupi_n_1445
    ^ csa_tree_add_48_2_groupi_n_1488));
 assign csa_tree_add_48_2_groupi_n_1621 = ((csa_tree_add_48_2_groupi_n_1513 & csa_tree_add_48_2_groupi_n_1559)
    | ((csa_tree_add_48_2_groupi_n_1559 & csa_tree_add_48_2_groupi_n_1489) | (csa_tree_add_48_2_groupi_n_1489
    & csa_tree_add_48_2_groupi_n_1513)));
 assign csa_tree_add_48_2_groupi_n_1622 = (csa_tree_add_48_2_groupi_n_1559 ^ (csa_tree_add_48_2_groupi_n_1489
    ^ csa_tree_add_48_2_groupi_n_1513));
 assign csa_tree_add_48_2_groupi_n_1620 = ~(csa_tree_add_48_2_groupi_n_1535 ^ csa_tree_add_48_2_groupi_n_1595);
 assign csa_tree_add_48_2_groupi_n_1619 = ~(csa_tree_add_48_2_groupi_n_1594 ^ csa_tree_add_48_2_groupi_n_1516);
 assign csa_tree_add_48_2_groupi_n_1625 = ~(csa_tree_add_48_2_groupi_n_1598 | csa_tree_add_48_2_groupi_n_96);
 assign csa_tree_add_48_2_groupi_n_1616 = ~(csa_tree_add_48_2_groupi_n_95 ^ csa_tree_add_48_2_groupi_n_1539);
 assign csa_tree_add_48_2_groupi_n_1618 = ~(csa_tree_add_48_2_groupi_n_97 & (csa_tree_add_48_2_groupi_n_1523
    | csa_tree_add_48_2_groupi_n_1590));
 assign csa_tree_add_48_2_groupi_n_1612 = (csa_tree_add_48_2_groupi_n_1575 & csa_tree_add_48_2_groupi_n_1534);
 assign csa_tree_add_48_2_groupi_n_1613 = (csa_tree_add_48_2_groupi_n_1575 ^ csa_tree_add_48_2_groupi_n_1534);
 assign csa_tree_add_48_2_groupi_n_1611 = ((csa_tree_add_48_2_groupi_n_1531 & csa_tree_add_48_2_groupi_n_1507)
    | ((csa_tree_add_48_2_groupi_n_1507 & csa_tree_add_48_2_groupi_n_1396) | (csa_tree_add_48_2_groupi_n_1396
    & csa_tree_add_48_2_groupi_n_1531)));
 assign csa_tree_add_48_2_groupi_n_1615 = (csa_tree_add_48_2_groupi_n_1507 ^ (csa_tree_add_48_2_groupi_n_1396
    ^ csa_tree_add_48_2_groupi_n_1531));
 assign csa_tree_add_48_2_groupi_n_1609 = ((csa_tree_add_48_2_groupi_n_1570 & csa_tree_add_48_2_groupi_n_1398)
    | ((csa_tree_add_48_2_groupi_n_1398 & csa_tree_add_48_2_groupi_n_1425) | (csa_tree_add_48_2_groupi_n_1425
    & csa_tree_add_48_2_groupi_n_1570)));
 assign csa_tree_add_48_2_groupi_n_1610 = (csa_tree_add_48_2_groupi_n_1398 ^ (csa_tree_add_48_2_groupi_n_1425
    ^ csa_tree_add_48_2_groupi_n_1570));
 assign csa_tree_add_48_2_groupi_n_1607 = ((csa_tree_add_48_2_groupi_n_1566 & csa_tree_add_48_2_groupi_n_1444)
    | ((csa_tree_add_48_2_groupi_n_1444 & csa_tree_add_48_2_groupi_n_1426) | (csa_tree_add_48_2_groupi_n_1426
    & csa_tree_add_48_2_groupi_n_1566)));
 assign csa_tree_add_48_2_groupi_n_1608 = (csa_tree_add_48_2_groupi_n_1444 ^ (csa_tree_add_48_2_groupi_n_1426
    ^ csa_tree_add_48_2_groupi_n_1566));
 assign csa_tree_add_48_2_groupi_n_1606 = (csa_tree_add_48_2_groupi_n_91 & csa_tree_add_48_2_groupi_n_1522);
 assign csa_tree_add_48_2_groupi_n_1614 = (csa_tree_add_48_2_groupi_n_91 ^ csa_tree_add_48_2_groupi_n_1522);
 assign csa_tree_add_48_2_groupi_n_1603 = ~(csa_tree_add_48_2_groupi_n_1535 | csa_tree_add_48_2_groupi_n_1595);
 assign csa_tree_add_48_2_groupi_n_1602 = ~(csa_tree_add_48_2_groupi_n_1594 | csa_tree_add_48_2_groupi_n_1516);
 assign csa_tree_add_48_2_groupi_n_1598 = ~(csa_tree_add_48_2_groupi_n_1548 | csa_tree_add_48_2_groupi_n_1543);
 assign csa_tree_add_48_2_groupi_n_1597 = (csa_tree_add_48_2_groupi_n_1535 & csa_tree_add_48_2_groupi_n_1595);
 assign csa_tree_add_48_2_groupi_n_1601 = (csa_tree_add_48_2_groupi_n_1579 ^ csa_tree_add_48_2_groupi_n_1413);
 assign csa_tree_add_48_2_groupi_n_1600 = ~(csa_tree_add_48_2_groupi_n_1525 & (csa_tree_add_48_2_groupi_n_1537
    | csa_tree_add_48_2_groupi_n_1528));
 assign csa_tree_add_48_2_groupi_n_1595 = ((csa_tree_add_48_2_groupi_n_1511 & csa_tree_add_48_2_groupi_n_1326)
    | ((csa_tree_add_48_2_groupi_n_1326 & csa_tree_add_48_2_groupi_n_1487) | (csa_tree_add_48_2_groupi_n_1487
    & csa_tree_add_48_2_groupi_n_1511)));
 assign csa_tree_add_48_2_groupi_n_1596 = (csa_tree_add_48_2_groupi_n_1326 ^ (csa_tree_add_48_2_groupi_n_1487
    ^ csa_tree_add_48_2_groupi_n_1511));
 assign csa_tree_add_48_2_groupi_n_1593 = ((csa_tree_add_48_2_groupi_n_1363 & csa_tree_add_48_2_groupi_n_1515)
    | ((csa_tree_add_48_2_groupi_n_1515 & csa_tree_add_48_2_groupi_n_65) | (csa_tree_add_48_2_groupi_n_65
    & csa_tree_add_48_2_groupi_n_1363)));
 assign csa_tree_add_48_2_groupi_n_1594 = (csa_tree_add_48_2_groupi_n_1515 ^ (csa_tree_add_48_2_groupi_n_65
    ^ csa_tree_add_48_2_groupi_n_1363));
 assign csa_tree_add_48_2_groupi_n_1590 = (csa_tree_add_48_2_groupi_n_87 & csa_tree_add_48_2_groupi_n_1536);
 assign csa_tree_add_48_2_groupi_n_1592 = (csa_tree_add_48_2_groupi_n_87 ^ csa_tree_add_48_2_groupi_n_1536);
 assign csa_tree_add_48_2_groupi_n_1589 = ((csa_tree_add_48_2_groupi_n_1529 & csa_tree_add_48_2_groupi_n_1400)
    | ((csa_tree_add_48_2_groupi_n_1400 & csa_tree_add_48_2_groupi_n_1485) | (csa_tree_add_48_2_groupi_n_1485
    & csa_tree_add_48_2_groupi_n_1529)));
 assign csa_tree_add_48_2_groupi_n_1591 = (csa_tree_add_48_2_groupi_n_1400 ^ (csa_tree_add_48_2_groupi_n_1485
    ^ csa_tree_add_48_2_groupi_n_1529));
 assign csa_tree_add_48_2_groupi_n_1584 = ~(csa_tree_add_48_2_groupi_n_1547 | (csa_tree_add_48_2_groupi_n_1546
    & csa_tree_add_48_2_groupi_n_1576));
 assign csa_tree_add_48_2_groupi_n_1582 = ((csa_tree_add_48_2_groupi_n_1399 & csa_tree_add_48_2_groupi_n_1465)
    | ((csa_tree_add_48_2_groupi_n_1465 & csa_tree_add_48_2_groupi_n_1484) | (csa_tree_add_48_2_groupi_n_1484
    & csa_tree_add_48_2_groupi_n_1399)));
 assign csa_tree_add_48_2_groupi_n_1583 = (csa_tree_add_48_2_groupi_n_1465 ^ (csa_tree_add_48_2_groupi_n_1484
    ^ csa_tree_add_48_2_groupi_n_1399));
 assign csa_tree_add_48_2_groupi_n_1581 = ~(csa_tree_add_48_2_groupi_n_91 | csa_tree_add_48_2_groupi_n_1522);
 assign csa_tree_add_48_2_groupi_n_1580 = ~(csa_tree_add_48_2_groupi_n_1574 & csa_tree_add_48_2_groupi_n_1533);
 assign csa_tree_add_48_2_groupi_n_1579 = ~((csa_tree_add_48_2_groupi_n_1518 & ~n_170) | (csa_tree_add_48_2_groupi_n_1538
    & n_170));
 assign csa_tree_add_48_2_groupi_n_1578 = ~(n_169 ^ csa_tree_add_48_2_groupi_n_1469);
 assign csa_tree_add_48_2_groupi_n_1577 = ~(csa_tree_add_48_2_groupi_n_1526 & (csa_tree_add_48_2_groupi_n_1527
    | csa_tree_add_48_2_groupi_n_1538));
 assign csa_tree_add_48_2_groupi_n_1576 = ~csa_tree_add_48_2_groupi_n_1517;
 assign csa_tree_add_48_2_groupi_n_1575 = ~csa_tree_add_48_2_groupi_n_1574;
 assign csa_tree_add_48_2_groupi_n_1572 = ((csa_tree_add_48_2_groupi_n_1446 & csa_tree_add_48_2_groupi_n_1424)
    | ((csa_tree_add_48_2_groupi_n_1424 & csa_tree_add_48_2_groupi_n_1230) | (csa_tree_add_48_2_groupi_n_1230
    & csa_tree_add_48_2_groupi_n_1446)));
 assign csa_tree_add_48_2_groupi_n_1573 = (csa_tree_add_48_2_groupi_n_1424 ^ (csa_tree_add_48_2_groupi_n_1230
    ^ csa_tree_add_48_2_groupi_n_1446));
 assign csa_tree_add_48_2_groupi_n_1570 = ((csa_tree_add_48_2_groupi_n_1459 & csa_tree_add_48_2_groupi_n_1165)
    | ((csa_tree_add_48_2_groupi_n_1165 & csa_tree_add_48_2_groupi_n_1337) | (csa_tree_add_48_2_groupi_n_1337
    & csa_tree_add_48_2_groupi_n_1459)));
 assign csa_tree_add_48_2_groupi_n_1571 = (csa_tree_add_48_2_groupi_n_1165 ^ (csa_tree_add_48_2_groupi_n_1337
    ^ csa_tree_add_48_2_groupi_n_1459));
 assign csa_tree_add_48_2_groupi_n_1566 = ((csa_tree_add_48_2_groupi_n_1466 & csa_tree_add_48_2_groupi_n_1375)
    | ((csa_tree_add_48_2_groupi_n_1375 & csa_tree_add_48_2_groupi_n_1460) | (csa_tree_add_48_2_groupi_n_1460
    & csa_tree_add_48_2_groupi_n_1466)));
 assign csa_tree_add_48_2_groupi_n_1567 = (csa_tree_add_48_2_groupi_n_1375 ^ (csa_tree_add_48_2_groupi_n_1460
    ^ csa_tree_add_48_2_groupi_n_1466));
 assign csa_tree_add_48_2_groupi_n_1564 = ((csa_tree_add_48_2_groupi_n_1442 & csa_tree_add_48_2_groupi_n_1447)
    | ((csa_tree_add_48_2_groupi_n_1447 & csa_tree_add_48_2_groupi_n_1225) | (csa_tree_add_48_2_groupi_n_1225
    & csa_tree_add_48_2_groupi_n_1442)));
 assign csa_tree_add_48_2_groupi_n_1565 = (csa_tree_add_48_2_groupi_n_1447 ^ (csa_tree_add_48_2_groupi_n_1225
    ^ csa_tree_add_48_2_groupi_n_1442));
 assign csa_tree_add_48_2_groupi_n_1560 = ((csa_tree_add_48_2_groupi_n_1436 & csa_tree_add_48_2_groupi_n_1443)
    | ((csa_tree_add_48_2_groupi_n_1443 & csa_tree_add_48_2_groupi_n_1208) | (csa_tree_add_48_2_groupi_n_1208
    & csa_tree_add_48_2_groupi_n_1436)));
 assign csa_tree_add_48_2_groupi_n_1561 = (csa_tree_add_48_2_groupi_n_1443 ^ (csa_tree_add_48_2_groupi_n_1208
    ^ csa_tree_add_48_2_groupi_n_1436));
 assign csa_tree_add_48_2_groupi_n_1558 = ((csa_tree_add_48_2_groupi_n_1464 & csa_tree_add_48_2_groupi_n_1467)
    | ((csa_tree_add_48_2_groupi_n_1467 & csa_tree_add_48_2_groupi_n_1438) | (csa_tree_add_48_2_groupi_n_1438
    & csa_tree_add_48_2_groupi_n_1464)));
 assign csa_tree_add_48_2_groupi_n_1559 = (csa_tree_add_48_2_groupi_n_1467 ^ (csa_tree_add_48_2_groupi_n_1438
    ^ csa_tree_add_48_2_groupi_n_1464));
 assign csa_tree_add_48_2_groupi_n_1557 = ((csa_tree_add_48_2_groupi_n_1404 & csa_tree_add_48_2_groupi_n_1437)
    | ((csa_tree_add_48_2_groupi_n_1437 & csa_tree_add_48_2_groupi_n_1264) | (csa_tree_add_48_2_groupi_n_1264
    & csa_tree_add_48_2_groupi_n_1404)));
 assign csa_tree_add_48_2_groupi_n_1574 = (csa_tree_add_48_2_groupi_n_1437 ^ (csa_tree_add_48_2_groupi_n_1264
    ^ csa_tree_add_48_2_groupi_n_1404));
 assign csa_tree_add_48_2_groupi_n_1548 = ~(n_169 | csa_tree_add_48_2_groupi_n_1469);
 assign csa_tree_add_48_2_groupi_n_1547 = ~(csa_tree_add_48_2_groupi_n_1540 | csa_tree_add_48_2_groupi_n_1498);
 assign csa_tree_add_48_2_groupi_n_1546 = ~(csa_tree_add_48_2_groupi_n_1540 & csa_tree_add_48_2_groupi_n_1498);
 assign csa_tree_add_48_2_groupi_n_1545 = ~(csa_tree_add_48_2_groupi_n_1532 | csa_tree_add_48_2_groupi_n_1519);
 assign csa_tree_add_48_2_groupi_n_1542 = ~(csa_tree_add_48_2_groupi_n_1532 & csa_tree_add_48_2_groupi_n_1519);
 assign csa_tree_add_48_2_groupi_n_1544 = ~((csa_tree_add_48_2_groupi_n_1455 & ~csa_tree_add_48_2_groupi_n_1520)
    | (csa_tree_add_48_2_groupi_n_1491 & csa_tree_add_48_2_groupi_n_1520));
 assign csa_tree_add_48_2_groupi_n_1541 = ~(csa_tree_add_48_2_groupi_n_1476 | (csa_tree_add_48_2_groupi_n_1482
    & csa_tree_add_48_2_groupi_n_1508));
 assign csa_tree_add_48_2_groupi_n_1543 = ~(csa_tree_add_48_2_groupi_n_1524 | csa_tree_add_48_2_groupi_n_90);
 assign csa_tree_add_48_2_groupi_n_1540 = ~csa_tree_add_48_2_groupi_n_1539;
 assign csa_tree_add_48_2_groupi_n_1538 = ~csa_tree_add_48_2_groupi_n_1518;
 assign csa_tree_add_48_2_groupi_n_1534 = ~csa_tree_add_48_2_groupi_n_1533;
 assign csa_tree_add_48_2_groupi_n_1532 = ~csa_tree_add_48_2_groupi_n_85;
 assign csa_tree_add_48_2_groupi_n_1531 = ((csa_tree_add_48_2_groupi_n_1368 & csa_tree_add_48_2_groupi_n_1461)
    | ((csa_tree_add_48_2_groupi_n_1461 & csa_tree_add_48_2_groupi_n_1354) | (csa_tree_add_48_2_groupi_n_1354
    & csa_tree_add_48_2_groupi_n_1368)));
 assign csa_tree_add_48_2_groupi_n_1539 = (csa_tree_add_48_2_groupi_n_1461 ^ (csa_tree_add_48_2_groupi_n_1354
    ^ csa_tree_add_48_2_groupi_n_1368));
 assign csa_tree_add_48_2_groupi_n_1536 = ((csa_tree_add_48_2_groupi_n_1364 & csa_tree_add_48_2_groupi_n_1361)
    | ((csa_tree_add_48_2_groupi_n_1361 & csa_tree_add_48_2_groupi_n_1381) | (csa_tree_add_48_2_groupi_n_1381
    & csa_tree_add_48_2_groupi_n_1364)));
 assign csa_tree_add_48_2_groupi_n_1537 = (csa_tree_add_48_2_groupi_n_1361 ^ (csa_tree_add_48_2_groupi_n_1381
    ^ csa_tree_add_48_2_groupi_n_1364));
 assign csa_tree_add_48_2_groupi_n_1533 = ((csa_tree_add_48_2_groupi_n_1486 & csa_tree_add_48_2_groupi_n_1405)
    | ((csa_tree_add_48_2_groupi_n_1405 & csa_tree_add_48_2_groupi_n_1371) | (csa_tree_add_48_2_groupi_n_1371
    & csa_tree_add_48_2_groupi_n_1486)));
 assign csa_tree_add_48_2_groupi_n_1535 = (csa_tree_add_48_2_groupi_n_1405 ^ (csa_tree_add_48_2_groupi_n_1371
    ^ csa_tree_add_48_2_groupi_n_1486));
 assign csa_tree_add_48_2_groupi_n_1529 = ((csa_tree_add_48_2_groupi_n_1422 & csa_tree_add_48_2_groupi_n_70)
    | ((csa_tree_add_48_2_groupi_n_70 & csa_tree_add_48_2_groupi_n_1402) | (csa_tree_add_48_2_groupi_n_1402
    & csa_tree_add_48_2_groupi_n_1422)));
 assign csa_tree_add_48_2_groupi_n_1530 = (csa_tree_add_48_2_groupi_n_70 ^ (csa_tree_add_48_2_groupi_n_1402
    ^ csa_tree_add_48_2_groupi_n_1422));
 assign csa_tree_add_48_2_groupi_n_1528 = ~(csa_tree_add_48_2_groupi_n_1520 | ~csa_tree_add_48_2_groupi_n_1455);
 assign csa_tree_add_48_2_groupi_n_1527 = ~(n_170 | csa_tree_add_48_2_groupi_n_1413);
 assign csa_tree_add_48_2_groupi_n_1526 = ~(n_170 & csa_tree_add_48_2_groupi_n_1413);
 assign csa_tree_add_48_2_groupi_n_1525 = ~(csa_tree_add_48_2_groupi_n_1491 & csa_tree_add_48_2_groupi_n_1520);
 assign csa_tree_add_48_2_groupi_n_1524 = ~(csa_tree_add_48_2_groupi_n_1477 | csa_tree_add_48_2_groupi_n_1499);
 assign csa_tree_add_48_2_groupi_n_1523 = (csa_tree_add_48_2_groupi_n_89 ^ csa_tree_add_48_2_groupi_n_1454);
 assign csa_tree_add_48_2_groupi_n_1521 = ~(csa_tree_add_48_2_groupi_n_1468 ^ (csa_tree_add_48_2_groupi_n_134
    ^ csa_tree_add_48_2_groupi_n_1360));
 assign csa_tree_add_48_2_groupi_n_1522 = ~(csa_tree_add_48_2_groupi_n_1502 & (csa_tree_add_48_2_groupi_n_1505
    | csa_tree_add_48_2_groupi_n_1471));
 assign csa_tree_add_48_2_groupi_n_1520 = ((csa_tree_add_48_2_groupi_n_1367 & n_173) | ((n_173 & csa_tree_add_48_2_groupi_n_46)
    | (csa_tree_add_48_2_groupi_n_46 & csa_tree_add_48_2_groupi_n_1367)));
 assign csa_tree_add_48_2_groupi_n_1515 = (n_173 ^ (csa_tree_add_48_2_groupi_n_46 ^ csa_tree_add_48_2_groupi_n_1367));
 assign csa_tree_add_48_2_groupi_n_1513 = ((csa_tree_add_48_2_groupi_n_1403 & csa_tree_add_48_2_groupi_n_1439)
    | ((csa_tree_add_48_2_groupi_n_1439 & csa_tree_add_48_2_groupi_n_1358) | (csa_tree_add_48_2_groupi_n_1358
    & csa_tree_add_48_2_groupi_n_1403)));
 assign csa_tree_add_48_2_groupi_n_1514 = (csa_tree_add_48_2_groupi_n_1439 ^ (csa_tree_add_48_2_groupi_n_1358
    ^ csa_tree_add_48_2_groupi_n_1403));
 assign csa_tree_add_48_2_groupi_n_1511 = ((csa_tree_add_48_2_groupi_n_1397 & csa_tree_add_48_2_groupi_n_1347)
    | ((csa_tree_add_48_2_groupi_n_1347 & csa_tree_add_48_2_groupi_n_1174) | (csa_tree_add_48_2_groupi_n_1174
    & csa_tree_add_48_2_groupi_n_1397)));
 assign csa_tree_add_48_2_groupi_n_1512 = (csa_tree_add_48_2_groupi_n_1347 ^ (csa_tree_add_48_2_groupi_n_1174
    ^ csa_tree_add_48_2_groupi_n_1397));
 assign csa_tree_add_48_2_groupi_n_1519 = ((csa_tree_add_48_2_groupi_n_1394 & csa_tree_add_48_2_groupi_n_1395)
    | ((csa_tree_add_48_2_groupi_n_1395 & csa_tree_add_48_2_groupi_n_1140) | (csa_tree_add_48_2_groupi_n_1140
    & csa_tree_add_48_2_groupi_n_1394)));
 assign csa_tree_add_48_2_groupi_n_1510 = (csa_tree_add_48_2_groupi_n_1395 ^ (csa_tree_add_48_2_groupi_n_1140
    ^ csa_tree_add_48_2_groupi_n_1394));
 assign csa_tree_add_48_2_groupi_n_1518 = ~(csa_tree_add_48_2_groupi_n_1506 & csa_tree_add_48_2_groupi_n_83);
 assign csa_tree_add_48_2_groupi_n_1517 = ~(csa_tree_add_48_2_groupi_n_1481 | (csa_tree_add_48_2_groupi_n_1480
    & csa_tree_add_48_2_groupi_n_1417));
 assign csa_tree_add_48_2_groupi_n_1516 = ~(csa_tree_add_48_2_groupi_n_86 & (csa_tree_add_48_2_groupi_n_1387
    | csa_tree_add_48_2_groupi_n_1483));
 assign csa_tree_add_48_2_groupi_n_1507 = ((csa_tree_add_48_2_groupi_n_1338 & csa_tree_add_48_2_groupi_n_1246)
    | ((csa_tree_add_48_2_groupi_n_1246 & csa_tree_add_48_2_groupi_n_1220) | (csa_tree_add_48_2_groupi_n_1220
    & csa_tree_add_48_2_groupi_n_1338)));
 assign csa_tree_add_48_2_groupi_n_1508 = (csa_tree_add_48_2_groupi_n_1246 ^ (csa_tree_add_48_2_groupi_n_1220
    ^ csa_tree_add_48_2_groupi_n_1338));
 assign csa_tree_add_48_2_groupi_n_1506 = ~(csa_tree_add_48_2_groupi_n_1421 & csa_tree_add_48_2_groupi_n_1366);
 assign csa_tree_add_48_2_groupi_n_1505 = ~(csa_tree_add_48_2_groupi_n_1454 | ~n_171);
 assign csa_tree_add_48_2_groupi_n_1502 = ~(csa_tree_add_48_2_groupi_n_1454 & ~n_171);
 assign csa_tree_add_48_2_groupi_n_1501 = ~((csa_tree_add_48_2_groupi_n_1418 & ~csa_tree_add_48_2_groupi_n_1451)
    | (csa_tree_add_48_2_groupi_n_1472 & csa_tree_add_48_2_groupi_n_1451));
 assign csa_tree_add_48_2_groupi_n_1500 = ~(csa_tree_add_48_2_groupi_n_1456 ^ csa_tree_add_48_2_groupi_n_1462);
 assign csa_tree_add_48_2_groupi_n_1495 = ~(csa_tree_add_48_2_groupi_n_1470 ^ csa_tree_add_48_2_groupi_n_75);
 assign csa_tree_add_48_2_groupi_n_1494 = ~((csa_tree_add_48_2_groupi_n_1412 & ~csa_tree_add_48_2_groupi_n_1415)
    | (csa_tree_add_48_2_groupi_n_1411 & csa_tree_add_48_2_groupi_n_1415));
 assign csa_tree_add_48_2_groupi_n_1499 = ~(csa_tree_add_48_2_groupi_n_1393 | (csa_tree_add_48_2_groupi_n_76
    & csa_tree_add_48_2_groupi_n_1452));
 assign csa_tree_add_48_2_groupi_n_1498 = ~(csa_tree_add_48_2_groupi_n_82 | csa_tree_add_48_2_groupi_n_1389);
 assign csa_tree_add_48_2_groupi_n_1493 = ~(csa_tree_add_48_2_groupi_n_1475 & csa_tree_add_48_2_groupi_n_1370);
 assign csa_tree_add_48_2_groupi_n_1492 = ~(csa_tree_add_48_2_groupi_n_1458 & (csa_tree_add_48_2_groupi_n_1457
    | csa_tree_add_48_2_groupi_n_1472));
 assign csa_tree_add_48_2_groupi_n_1491 = ~csa_tree_add_48_2_groupi_n_1455;
 assign csa_tree_add_48_2_groupi_n_1488 = ((csa_tree_add_48_2_groupi_n_1357 & csa_tree_add_48_2_groupi_n_1376)
    | ((csa_tree_add_48_2_groupi_n_1376 & csa_tree_add_48_2_groupi_n_1162) | (csa_tree_add_48_2_groupi_n_1162
    & csa_tree_add_48_2_groupi_n_1357)));
 assign csa_tree_add_48_2_groupi_n_1489 = (csa_tree_add_48_2_groupi_n_1376 ^ (csa_tree_add_48_2_groupi_n_1162
    ^ csa_tree_add_48_2_groupi_n_1357));
 assign csa_tree_add_48_2_groupi_n_1486 = ((csa_tree_add_48_2_groupi_n_1173 & csa_tree_add_48_2_groupi_n_1372)
    | ((csa_tree_add_48_2_groupi_n_1372 & csa_tree_add_48_2_groupi_n_1248) | (csa_tree_add_48_2_groupi_n_1248
    & csa_tree_add_48_2_groupi_n_1173)));
 assign csa_tree_add_48_2_groupi_n_1487 = (csa_tree_add_48_2_groupi_n_1372 ^ (csa_tree_add_48_2_groupi_n_1248
    ^ csa_tree_add_48_2_groupi_n_1173));
 assign csa_tree_add_48_2_groupi_n_1484 = ((csa_tree_add_48_2_groupi_n_1401 & csa_tree_add_48_2_groupi_n_1172)
    | ((csa_tree_add_48_2_groupi_n_1172 & csa_tree_add_48_2_groupi_n_1170) | (csa_tree_add_48_2_groupi_n_1170
    & csa_tree_add_48_2_groupi_n_1401)));
 assign csa_tree_add_48_2_groupi_n_1485 = (csa_tree_add_48_2_groupi_n_1172 ^ (csa_tree_add_48_2_groupi_n_1170
    ^ csa_tree_add_48_2_groupi_n_1401));
 assign csa_tree_add_48_2_groupi_n_1483 = (csa_tree_add_48_2_groupi_n_72 & csa_tree_add_48_2_groupi_n_1378);
 assign csa_tree_add_48_2_groupi_n_1490 = (csa_tree_add_48_2_groupi_n_72 ^ csa_tree_add_48_2_groupi_n_1378);
 assign csa_tree_add_48_2_groupi_n_1482 = ~(csa_tree_add_48_2_groupi_n_1415 & csa_tree_add_48_2_groupi_n_1412);
 assign csa_tree_add_48_2_groupi_n_1481 = ~(csa_tree_add_48_2_groupi_n_1414 | n_172);
 assign csa_tree_add_48_2_groupi_n_1480 = ~(csa_tree_add_48_2_groupi_n_1414 & n_172);
 assign csa_tree_add_48_2_groupi_n_1477 = ~(csa_tree_add_48_2_groupi_n_1470 | csa_tree_add_48_2_groupi_n_75);
 assign csa_tree_add_48_2_groupi_n_1476 = ~(csa_tree_add_48_2_groupi_n_1415 | csa_tree_add_48_2_groupi_n_1412);
 assign csa_tree_add_48_2_groupi_n_1475 = ~(csa_tree_add_48_2_groupi_n_1468 & csa_tree_add_48_2_groupi_n_61);
 assign csa_tree_add_48_2_groupi_n_1474 = ~((csa_tree_add_48_2_groupi_n_1365 & ~csa_tree_add_48_2_groupi_n_1386)
    | (csa_tree_add_48_2_groupi_n_1407 & csa_tree_add_48_2_groupi_n_1386));
 assign csa_tree_add_48_2_groupi_n_1473 = ~(csa_tree_add_48_2_groupi_n_1420 & (csa_tree_add_48_2_groupi_n_1419
    | csa_tree_add_48_2_groupi_n_1386));
 assign csa_tree_add_48_2_groupi_n_1472 = ~csa_tree_add_48_2_groupi_n_1418;
 assign csa_tree_add_48_2_groupi_n_1471 = ~csa_tree_add_48_2_groupi_n_79;
 assign csa_tree_add_48_2_groupi_n_1466 = ((csa_tree_add_48_2_groupi_n_1164 & csa_tree_add_48_2_groupi_n_1286)
    | ((csa_tree_add_48_2_groupi_n_1286 & csa_tree_add_48_2_groupi_n_1295) | (csa_tree_add_48_2_groupi_n_1295
    & csa_tree_add_48_2_groupi_n_1164)));
 assign csa_tree_add_48_2_groupi_n_1467 = (csa_tree_add_48_2_groupi_n_1286 ^ (csa_tree_add_48_2_groupi_n_1295
    ^ csa_tree_add_48_2_groupi_n_1164));
 assign csa_tree_add_48_2_groupi_n_1469 = ((csa_tree_add_48_2_groupi_n_1339 & csa_tree_add_48_2_groupi_n_53)
    | ((csa_tree_add_48_2_groupi_n_53 & csa_tree_add_48_2_groupi_n_1185) | (csa_tree_add_48_2_groupi_n_1185
    & csa_tree_add_48_2_groupi_n_1339)));
 assign csa_tree_add_48_2_groupi_n_1470 = (csa_tree_add_48_2_groupi_n_53 ^ (csa_tree_add_48_2_groupi_n_1185
    ^ csa_tree_add_48_2_groupi_n_1339));
 assign csa_tree_add_48_2_groupi_n_1464 = ((csa_tree_add_48_2_groupi_n_1169 & csa_tree_add_48_2_groupi_n_1178)
    | ((csa_tree_add_48_2_groupi_n_1178 & csa_tree_add_48_2_groupi_n_1296) | (csa_tree_add_48_2_groupi_n_1296
    & csa_tree_add_48_2_groupi_n_1169)));
 assign csa_tree_add_48_2_groupi_n_1465 = (csa_tree_add_48_2_groupi_n_1178 ^ (csa_tree_add_48_2_groupi_n_1296
    ^ csa_tree_add_48_2_groupi_n_1169));
 assign csa_tree_add_48_2_groupi_n_1462 = ((csa_tree_add_48_2_groupi_n_1257 & csa_tree_add_48_2_groupi_n_1298)
    | ((csa_tree_add_48_2_groupi_n_1298 & csa_tree_add_48_2_groupi_n_1243) | (csa_tree_add_48_2_groupi_n_1243
    & csa_tree_add_48_2_groupi_n_1257)));
 assign csa_tree_add_48_2_groupi_n_1463 = (csa_tree_add_48_2_groupi_n_1298 ^ (csa_tree_add_48_2_groupi_n_1243
    ^ csa_tree_add_48_2_groupi_n_1257));
 assign csa_tree_add_48_2_groupi_n_1468 = ((csa_tree_add_48_2_groupi_n_1287 & csa_tree_add_48_2_groupi_n_1289)
    | ((csa_tree_add_48_2_groupi_n_1289 & csa_tree_add_48_2_groupi_n_1213) | (csa_tree_add_48_2_groupi_n_1213
    & csa_tree_add_48_2_groupi_n_1287)));
 assign csa_tree_add_48_2_groupi_n_1461 = (csa_tree_add_48_2_groupi_n_1289 ^ (csa_tree_add_48_2_groupi_n_1213
    ^ csa_tree_add_48_2_groupi_n_1287));
 assign csa_tree_add_48_2_groupi_n_1459 = ((csa_tree_add_48_2_groupi_n_1161 & csa_tree_add_48_2_groupi_n_1163)
    | ((csa_tree_add_48_2_groupi_n_1163 & csa_tree_add_48_2_groupi_n_1285) | (csa_tree_add_48_2_groupi_n_1285
    & csa_tree_add_48_2_groupi_n_1161)));
 assign csa_tree_add_48_2_groupi_n_1460 = (csa_tree_add_48_2_groupi_n_1163 ^ (csa_tree_add_48_2_groupi_n_1285
    ^ csa_tree_add_48_2_groupi_n_1161));
 assign csa_tree_add_48_2_groupi_n_1458 = ~(csa_tree_add_48_2_groupi_n_1451 & csa_tree_add_48_2_groupi_n_1406);
 assign csa_tree_add_48_2_groupi_n_1457 = ~(csa_tree_add_48_2_groupi_n_1451 | csa_tree_add_48_2_groupi_n_1406);
 assign csa_tree_add_48_2_groupi_n_1456 = ~(csa_tree_add_48_2_groupi_n_1383 ^ csa_tree_add_48_2_groupi_n_1179);
 assign csa_tree_add_48_2_groupi_n_1453 = ~((csa_tree_add_48_2_groupi_n_1410 & ~n_175) | (csa_tree_add_48_2_groupi_n_1377
    & n_175));
 assign csa_tree_add_48_2_groupi_n_1455 = (csa_tree_add_48_2_groupi_n_77 ^ csa_tree_add_48_2_groupi_n_1379);
 assign csa_tree_add_48_2_groupi_n_1454 = ~(csa_tree_add_48_2_groupi_n_1318 & (csa_tree_add_48_2_groupi_n_1324
    | csa_tree_add_48_2_groupi_n_1409));
 assign csa_tree_add_48_2_groupi_n_1448 = ((csa_tree_add_48_2_groupi_n_1211 & csa_tree_add_48_2_groupi_n_1250)
    | ((csa_tree_add_48_2_groupi_n_1250 & csa_tree_add_48_2_groupi_n_1217) | (csa_tree_add_48_2_groupi_n_1217
    & csa_tree_add_48_2_groupi_n_1211)));
 assign csa_tree_add_48_2_groupi_n_1449 = (csa_tree_add_48_2_groupi_n_1250 ^ (csa_tree_add_48_2_groupi_n_1217
    ^ csa_tree_add_48_2_groupi_n_1211));
 assign csa_tree_add_48_2_groupi_n_1446 = ((csa_tree_add_48_2_groupi_n_1207 & csa_tree_add_48_2_groupi_n_1227)
    | ((csa_tree_add_48_2_groupi_n_1227 & csa_tree_add_48_2_groupi_n_1209) | (csa_tree_add_48_2_groupi_n_1209
    & csa_tree_add_48_2_groupi_n_1207)));
 assign csa_tree_add_48_2_groupi_n_1447 = (csa_tree_add_48_2_groupi_n_1227 ^ (csa_tree_add_48_2_groupi_n_1209
    ^ csa_tree_add_48_2_groupi_n_1207));
 assign csa_tree_add_48_2_groupi_n_1444 = ((csa_tree_add_48_2_groupi_n_1168 & csa_tree_add_48_2_groupi_n_1291)
    | ((csa_tree_add_48_2_groupi_n_1291 & csa_tree_add_48_2_groupi_n_1166) | (csa_tree_add_48_2_groupi_n_1166
    & csa_tree_add_48_2_groupi_n_1168)));
 assign csa_tree_add_48_2_groupi_n_1445 = (csa_tree_add_48_2_groupi_n_1291 ^ (csa_tree_add_48_2_groupi_n_1166
    ^ csa_tree_add_48_2_groupi_n_1168));
 assign csa_tree_add_48_2_groupi_n_1442 = ((csa_tree_add_48_2_groupi_n_1263 & csa_tree_add_48_2_groupi_n_1210)
    | ((csa_tree_add_48_2_groupi_n_1210 & csa_tree_add_48_2_groupi_n_1265) | (csa_tree_add_48_2_groupi_n_1265
    & csa_tree_add_48_2_groupi_n_1263)));
 assign csa_tree_add_48_2_groupi_n_1443 = (csa_tree_add_48_2_groupi_n_1210 ^ (csa_tree_add_48_2_groupi_n_1265
    ^ csa_tree_add_48_2_groupi_n_1263));
 assign csa_tree_add_48_2_groupi_n_1440 = ((csa_tree_add_48_2_groupi_n_1253 & csa_tree_add_48_2_groupi_n_1218)
    | ((csa_tree_add_48_2_groupi_n_1218 & csa_tree_add_48_2_groupi_n_1259) | (csa_tree_add_48_2_groupi_n_1259
    & csa_tree_add_48_2_groupi_n_1253)));
 assign csa_tree_add_48_2_groupi_n_1441 = (csa_tree_add_48_2_groupi_n_1218 ^ (csa_tree_add_48_2_groupi_n_1259
    ^ csa_tree_add_48_2_groupi_n_1253));
 assign csa_tree_add_48_2_groupi_n_1438 = ((csa_tree_add_48_2_groupi_n_1292 & csa_tree_add_48_2_groupi_n_1176)
    | ((csa_tree_add_48_2_groupi_n_1176 & csa_tree_add_48_2_groupi_n_1171) | (csa_tree_add_48_2_groupi_n_1171
    & csa_tree_add_48_2_groupi_n_1292)));
 assign csa_tree_add_48_2_groupi_n_1439 = (csa_tree_add_48_2_groupi_n_1176 ^ (csa_tree_add_48_2_groupi_n_1171
    ^ csa_tree_add_48_2_groupi_n_1292));
 assign csa_tree_add_48_2_groupi_n_1436 = ((csa_tree_add_48_2_groupi_n_1251 & csa_tree_add_48_2_groupi_n_1266)
    | ((csa_tree_add_48_2_groupi_n_1266 & csa_tree_add_48_2_groupi_n_1238) | (csa_tree_add_48_2_groupi_n_1238
    & csa_tree_add_48_2_groupi_n_1251)));
 assign csa_tree_add_48_2_groupi_n_1437 = (csa_tree_add_48_2_groupi_n_1266 ^ (csa_tree_add_48_2_groupi_n_1238
    ^ csa_tree_add_48_2_groupi_n_1251));
 assign csa_tree_add_48_2_groupi_n_1433 = ((csa_tree_add_48_2_groupi_n_1229 & csa_tree_add_48_2_groupi_n_1260)
    | ((csa_tree_add_48_2_groupi_n_1260 & csa_tree_add_48_2_groupi_n_1240) | (csa_tree_add_48_2_groupi_n_1240
    & csa_tree_add_48_2_groupi_n_1229)));
 assign csa_tree_add_48_2_groupi_n_1434 = (csa_tree_add_48_2_groupi_n_1260 ^ (csa_tree_add_48_2_groupi_n_1240
    ^ csa_tree_add_48_2_groupi_n_1229));
 assign csa_tree_add_48_2_groupi_n_1431 = ((csa_tree_add_48_2_groupi_n_1234 & csa_tree_add_48_2_groupi_n_1232)
    | ((csa_tree_add_48_2_groupi_n_1232 & csa_tree_add_48_2_groupi_n_1249) | (csa_tree_add_48_2_groupi_n_1249
    & csa_tree_add_48_2_groupi_n_1234)));
 assign csa_tree_add_48_2_groupi_n_1432 = (csa_tree_add_48_2_groupi_n_1232 ^ (csa_tree_add_48_2_groupi_n_1249
    ^ csa_tree_add_48_2_groupi_n_1234));
 assign csa_tree_add_48_2_groupi_n_1429 = ((csa_tree_add_48_2_groupi_n_1261 & csa_tree_add_48_2_groupi_n_1244)
    | ((csa_tree_add_48_2_groupi_n_1244 & csa_tree_add_48_2_groupi_n_1231) | (csa_tree_add_48_2_groupi_n_1231
    & csa_tree_add_48_2_groupi_n_1261)));
 assign csa_tree_add_48_2_groupi_n_1430 = (csa_tree_add_48_2_groupi_n_1244 ^ (csa_tree_add_48_2_groupi_n_1231
    ^ csa_tree_add_48_2_groupi_n_1261));
 assign csa_tree_add_48_2_groupi_n_1427 = ((csa_tree_add_48_2_groupi_n_1336 & csa_tree_add_48_2_groupi_n_1228)
    | ((csa_tree_add_48_2_groupi_n_1228 & csa_tree_add_48_2_groupi_n_876) | (csa_tree_add_48_2_groupi_n_876
    & csa_tree_add_48_2_groupi_n_1336)));
 assign csa_tree_add_48_2_groupi_n_1428 = (csa_tree_add_48_2_groupi_n_1228 ^ (csa_tree_add_48_2_groupi_n_876
    ^ csa_tree_add_48_2_groupi_n_1336));
 assign csa_tree_add_48_2_groupi_n_1425 = ((csa_tree_add_48_2_groupi_n_1290 & csa_tree_add_48_2_groupi_n_1222)
    | ((csa_tree_add_48_2_groupi_n_1222 & csa_tree_add_48_2_groupi_n_1121) | (csa_tree_add_48_2_groupi_n_1121
    & csa_tree_add_48_2_groupi_n_1290)));
 assign csa_tree_add_48_2_groupi_n_1426 = (csa_tree_add_48_2_groupi_n_1222 ^ (csa_tree_add_48_2_groupi_n_1121
    ^ csa_tree_add_48_2_groupi_n_1290));
 assign csa_tree_add_48_2_groupi_n_1423 = ((csa_tree_add_48_2_groupi_n_1224 & csa_tree_add_48_2_groupi_n_1241)
    | ((csa_tree_add_48_2_groupi_n_1241 & csa_tree_add_48_2_groupi_n_1226) | (csa_tree_add_48_2_groupi_n_1226
    & csa_tree_add_48_2_groupi_n_1224)));
 assign csa_tree_add_48_2_groupi_n_1424 = (csa_tree_add_48_2_groupi_n_1241 ^ (csa_tree_add_48_2_groupi_n_1226
    ^ csa_tree_add_48_2_groupi_n_1224));
 assign csa_tree_add_48_2_groupi_n_1422 = ((csa_tree_add_48_2_groupi_n_1245 & csa_tree_add_48_2_groupi_n_1132)
    | ((csa_tree_add_48_2_groupi_n_1132 & csa_tree_add_48_2_groupi_n_1186) | (csa_tree_add_48_2_groupi_n_1186
    & csa_tree_add_48_2_groupi_n_1245)));
 assign csa_tree_add_48_2_groupi_n_1451 = (csa_tree_add_48_2_groupi_n_1132 ^ (csa_tree_add_48_2_groupi_n_1186
    ^ csa_tree_add_48_2_groupi_n_1245));
 assign csa_tree_add_48_2_groupi_n_1421 = ~(n_175 & csa_tree_add_48_2_groupi_n_1410);
 assign csa_tree_add_48_2_groupi_n_1420 = ~(csa_tree_add_48_2_groupi_n_1408 & csa_tree_add_48_2_groupi_n_1407);
 assign csa_tree_add_48_2_groupi_n_1419 = ~(csa_tree_add_48_2_groupi_n_1408 | csa_tree_add_48_2_groupi_n_1407);
 assign csa_tree_add_48_2_groupi_n_1450 = ~(csa_tree_add_48_2_groupi_n_1390 | csa_tree_add_48_2_groupi_n_1391);
 assign csa_tree_add_48_2_groupi_n_1418 = ~(csa_tree_add_48_2_groupi_n_1384 & csa_tree_add_48_2_groupi_n_1320);
 assign csa_tree_add_48_2_groupi_n_1417 = ~(csa_tree_add_48_2_groupi_n_1319 & (csa_tree_add_48_2_groupi_n_1280
    | csa_tree_add_48_2_groupi_n_1328));
 assign csa_tree_add_48_2_groupi_n_1415 = ~(csa_tree_add_48_2_groupi_n_1388 | (csa_tree_add_48_2_groupi_n_1346
    & csa_tree_add_48_2_groupi_n_1271));
 assign csa_tree_add_48_2_groupi_n_1414 = ~(csa_tree_add_48_2_groupi_n_1373 | (csa_tree_add_48_2_groupi_n_78
    & csa_tree_add_48_2_groupi_n_1316));
 assign csa_tree_add_48_2_groupi_n_1412 = ~csa_tree_add_48_2_groupi_n_1411;
 assign csa_tree_add_48_2_groupi_n_1410 = ~csa_tree_add_48_2_groupi_n_1377;
 assign csa_tree_add_48_2_groupi_n_1409 = ~csa_tree_add_48_2_groupi_n_1379;
 assign csa_tree_add_48_2_groupi_n_1407 = ~csa_tree_add_48_2_groupi_n_1365;
 assign csa_tree_add_48_2_groupi_n_1411 = ((csa_tree_add_48_2_groupi_n_1216 & csa_tree_add_48_2_groupi_n_1288)
    | ((csa_tree_add_48_2_groupi_n_1288 & csa_tree_add_48_2_groupi_n_1214) | (csa_tree_add_48_2_groupi_n_1214
    & csa_tree_add_48_2_groupi_n_1216)));
 assign csa_tree_add_48_2_groupi_n_1413 = (csa_tree_add_48_2_groupi_n_1288 ^ (csa_tree_add_48_2_groupi_n_1214
    ^ csa_tree_add_48_2_groupi_n_1216));
 assign csa_tree_add_48_2_groupi_n_1404 = ((csa_tree_add_48_2_groupi_n_1247 & csa_tree_add_48_2_groupi_n_1239)
    | ((csa_tree_add_48_2_groupi_n_1239 & csa_tree_add_48_2_groupi_n_1252) | (csa_tree_add_48_2_groupi_n_1252
    & csa_tree_add_48_2_groupi_n_1247)));
 assign csa_tree_add_48_2_groupi_n_1405 = (csa_tree_add_48_2_groupi_n_1239 ^ (csa_tree_add_48_2_groupi_n_1252
    ^ csa_tree_add_48_2_groupi_n_1247));
 assign csa_tree_add_48_2_groupi_n_1403 = ((csa_tree_add_48_2_groupi_n_1267 & csa_tree_add_48_2_groupi_n_1242)
    | ((csa_tree_add_48_2_groupi_n_1242 & csa_tree_add_48_2_groupi_n_1198) | (csa_tree_add_48_2_groupi_n_1198
    & csa_tree_add_48_2_groupi_n_1267)));
 assign csa_tree_add_48_2_groupi_n_1408 = (csa_tree_add_48_2_groupi_n_1242 ^ (csa_tree_add_48_2_groupi_n_1198
    ^ csa_tree_add_48_2_groupi_n_1267));
 assign csa_tree_add_48_2_groupi_n_1401 = ((csa_tree_add_48_2_groupi_n_1236 & csa_tree_add_48_2_groupi_n_1088)
    | ((csa_tree_add_48_2_groupi_n_1088 & csa_tree_add_48_2_groupi_n_918) | (csa_tree_add_48_2_groupi_n_918
    & csa_tree_add_48_2_groupi_n_1236)));
 assign csa_tree_add_48_2_groupi_n_1402 = (csa_tree_add_48_2_groupi_n_1088 ^ (csa_tree_add_48_2_groupi_n_918
    ^ csa_tree_add_48_2_groupi_n_1236));
 assign csa_tree_add_48_2_groupi_n_1399 = ((csa_tree_add_48_2_groupi_n_1256 & csa_tree_add_48_2_groupi_n_1293)
    | ((csa_tree_add_48_2_groupi_n_1293 & csa_tree_add_48_2_groupi_n_1233) | (csa_tree_add_48_2_groupi_n_1233
    & csa_tree_add_48_2_groupi_n_1256)));
 assign csa_tree_add_48_2_groupi_n_1400 = (csa_tree_add_48_2_groupi_n_1293 ^ (csa_tree_add_48_2_groupi_n_1233
    ^ csa_tree_add_48_2_groupi_n_1256));
 assign csa_tree_add_48_2_groupi_n_1397 = ((csa_tree_add_48_2_groupi_n_1221 & csa_tree_add_48_2_groupi_n_920)
    | ((csa_tree_add_48_2_groupi_n_920 & csa_tree_add_48_2_groupi_n_1120) | (csa_tree_add_48_2_groupi_n_1120
    & csa_tree_add_48_2_groupi_n_1221)));
 assign csa_tree_add_48_2_groupi_n_1398 = (csa_tree_add_48_2_groupi_n_920 ^ (csa_tree_add_48_2_groupi_n_1120
    ^ csa_tree_add_48_2_groupi_n_1221));
 assign csa_tree_add_48_2_groupi_n_1395 = ((csa_tree_add_48_2_groupi_n_1237 & csa_tree_add_48_2_groupi_n_1141)
    | ((csa_tree_add_48_2_groupi_n_1141 & csa_tree_add_48_2_groupi_n_1087) | (csa_tree_add_48_2_groupi_n_1087
    & csa_tree_add_48_2_groupi_n_1237)));
 assign csa_tree_add_48_2_groupi_n_1396 = (csa_tree_add_48_2_groupi_n_1141 ^ (csa_tree_add_48_2_groupi_n_1087
    ^ csa_tree_add_48_2_groupi_n_1237));
 assign csa_tree_add_48_2_groupi_n_1394 = ((csa_tree_add_48_2_groupi_n_1219 & csa_tree_add_48_2_groupi_n_1223)
    | ((csa_tree_add_48_2_groupi_n_1223 & csa_tree_add_48_2_groupi_n_1090) | (csa_tree_add_48_2_groupi_n_1090
    & csa_tree_add_48_2_groupi_n_1219)));
 assign csa_tree_add_48_2_groupi_n_1406 = (csa_tree_add_48_2_groupi_n_1223 ^ (csa_tree_add_48_2_groupi_n_1090
    ^ csa_tree_add_48_2_groupi_n_1219));
 assign csa_tree_add_48_2_groupi_n_1393 = ~(n_174 | ~csa_tree_add_48_2_groupi_n_1311);
 assign csa_tree_add_48_2_groupi_n_1392 = ~(csa_tree_add_48_2_groupi_n_1380 | csa_tree_add_48_2_groupi_n_1302);
 assign csa_tree_add_48_2_groupi_n_1391 = ~(n_176 | csa_tree_add_48_2_groupi_n_1302);
 assign csa_tree_add_48_2_groupi_n_1390 = ~(csa_tree_add_48_2_groupi_n_1380 | csa_tree_add_48_2_groupi_n_1301);
 assign csa_tree_add_48_2_groupi_n_1389 = ~(n_176 | csa_tree_add_48_2_groupi_n_1301);
 assign csa_tree_add_48_2_groupi_n_1388 = ~(csa_tree_add_48_2_groupi_n_1346 | csa_tree_add_48_2_groupi_n_1271);
 assign csa_tree_add_48_2_groupi_n_1384 = ~(csa_tree_add_48_2_groupi_n_1335 & csa_tree_add_48_2_groupi_n_1271);
 assign csa_tree_add_48_2_groupi_n_1383 = ~(csa_tree_add_48_2_groupi_n_1348 ^ csa_tree_add_48_2_groupi_n_1133);
 assign csa_tree_add_48_2_groupi_n_1387 = (csa_tree_add_48_2_groupi_n_1341 ^ csa_tree_add_48_2_groupi_n_38);
 assign csa_tree_add_48_2_groupi_n_1382 = (csa_tree_add_48_2_groupi_n_1356 ^ csa_tree_add_48_2_groupi_n_1281);
 assign csa_tree_add_48_2_groupi_n_1386 = ~(csa_tree_add_48_2_groupi_n_1355 | (csa_tree_add_48_2_groupi_n_64
    & csa_tree_add_48_2_groupi_n_1281));
 assign csa_tree_add_48_2_groupi_n_1381 = (csa_tree_add_48_2_groupi_n_74 ^ csa_tree_add_48_2_groupi_n_1189);
 assign csa_tree_add_48_2_groupi_n_1380 = ~n_176;
 assign csa_tree_add_48_2_groupi_n_1375 = ((csa_tree_add_48_2_groupi_n_1177 & csa_tree_add_48_2_groupi_n_916)
    | ((csa_tree_add_48_2_groupi_n_916 & csa_tree_add_48_2_groupi_n_1175) | (csa_tree_add_48_2_groupi_n_1175
    & csa_tree_add_48_2_groupi_n_1177)));
 assign csa_tree_add_48_2_groupi_n_1376 = (csa_tree_add_48_2_groupi_n_916 ^ (csa_tree_add_48_2_groupi_n_1175
    ^ csa_tree_add_48_2_groupi_n_1177));
 assign csa_tree_add_48_2_groupi_n_1373 = (csa_tree_add_48_2_groupi_n_37 & csa_tree_add_48_2_groupi_n_1191);
 assign csa_tree_add_48_2_groupi_n_1374 = (csa_tree_add_48_2_groupi_n_37 ^ csa_tree_add_48_2_groupi_n_1191);
 assign csa_tree_add_48_2_groupi_n_1371 = ((csa_tree_add_48_2_groupi_n_1294 & csa_tree_add_48_2_groupi_n_914)
    | ((csa_tree_add_48_2_groupi_n_914 & csa_tree_add_48_2_groupi_n_1038) | (csa_tree_add_48_2_groupi_n_1038
    & csa_tree_add_48_2_groupi_n_1294)));
 assign csa_tree_add_48_2_groupi_n_1372 = (csa_tree_add_48_2_groupi_n_914 ^ (csa_tree_add_48_2_groupi_n_1038
    ^ csa_tree_add_48_2_groupi_n_1294));
 assign csa_tree_add_48_2_groupi_n_1370 = ~(csa_tree_add_48_2_groupi_n_134 & csa_tree_add_48_2_groupi_n_1360);
 assign csa_tree_add_48_2_groupi_n_1368 = ~(csa_tree_add_48_2_groupi_n_1334 & (csa_tree_add_48_2_groupi_n_1333
    | csa_tree_add_48_2_groupi_n_1277));
 assign csa_tree_add_48_2_groupi_n_1379 = ~(csa_tree_add_48_2_groupi_n_1206 & (csa_tree_add_48_2_groupi_n_1200
    | csa_tree_add_48_2_groupi_n_1307));
 assign csa_tree_add_48_2_groupi_n_1367 = ~(csa_tree_add_48_2_groupi_n_1201 & (csa_tree_add_48_2_groupi_n_1193
    | csa_tree_add_48_2_groupi_n_1205));
 assign csa_tree_add_48_2_groupi_n_1378 = ~(csa_tree_add_48_2_groupi_n_1199 | (csa_tree_add_48_2_groupi_n_1204
    & csa_tree_add_48_2_groupi_n_1310));
 assign csa_tree_add_48_2_groupi_n_1377 = ~(csa_tree_add_48_2_groupi_n_1350 & csa_tree_add_48_2_groupi_n_1202);
 assign csa_tree_add_48_2_groupi_n_1364 = ~(csa_tree_add_48_2_groupi_n_1323 | (csa_tree_add_48_2_groupi_n_1322
    & csa_tree_add_48_2_groupi_n_1305));
 assign csa_tree_add_48_2_groupi_n_1363 = ~(csa_tree_add_48_2_groupi_n_1352 & csa_tree_add_48_2_groupi_n_73);
 assign csa_tree_add_48_2_groupi_n_1366 = ~(csa_tree_add_48_2_groupi_n_1351 & csa_tree_add_48_2_groupi_n_1321);
 assign csa_tree_add_48_2_groupi_n_1365 = ~(csa_tree_add_48_2_groupi_n_1353 | csa_tree_add_48_2_groupi_n_1203);
 assign csa_tree_add_48_2_groupi_n_1361 = ~(csa_tree_add_48_2_groupi_n_1282 ^ csa_tree_add_48_2_groupi_n_1194);
 assign csa_tree_add_48_2_groupi_n_1357 = ((csa_tree_add_48_2_groupi_n_1255 & csa_tree_add_48_2_groupi_n_915)
    | ((csa_tree_add_48_2_groupi_n_915 & csa_tree_add_48_2_groupi_n_947) | (csa_tree_add_48_2_groupi_n_947
    & csa_tree_add_48_2_groupi_n_1255)));
 assign csa_tree_add_48_2_groupi_n_1358 = (csa_tree_add_48_2_groupi_n_915 ^ (csa_tree_add_48_2_groupi_n_947
    ^ csa_tree_add_48_2_groupi_n_1255));
 assign csa_tree_add_48_2_groupi_n_1355 = (csa_tree_add_48_2_groupi_n_1273 & csa_tree_add_48_2_groupi_n_1274);
 assign csa_tree_add_48_2_groupi_n_1356 = (csa_tree_add_48_2_groupi_n_1273 ^ csa_tree_add_48_2_groupi_n_1274);
 assign csa_tree_add_48_2_groupi_n_1360 = (csa_tree_add_48_2_groupi_n_1215 & csa_tree_add_48_2_groupi_n_1122);
 assign csa_tree_add_48_2_groupi_n_1354 = (csa_tree_add_48_2_groupi_n_1215 ^ csa_tree_add_48_2_groupi_n_1122);
 assign csa_tree_add_48_2_groupi_n_1353 = ~(csa_tree_add_48_2_groupi_n_1197 | csa_tree_add_48_2_groupi_n_60);
 assign csa_tree_add_48_2_groupi_n_1352 = ~(csa_tree_add_48_2_groupi_n_71 & csa_tree_add_48_2_groupi_n_1303);
 assign csa_tree_add_48_2_groupi_n_1351 = ~(csa_tree_add_48_2_groupi_n_1152 & (csa_tree_add_48_2_groupi_n_1189
    | csa_tree_add_48_2_groupi_n_1268));
 assign csa_tree_add_48_2_groupi_n_1350 = ~(csa_tree_add_48_2_groupi_n_1309 & (csa_tree_add_48_2_groupi_n_1131
    | csa_tree_add_48_2_groupi_n_1182));
 assign csa_tree_add_48_2_groupi_n_1349 = ~((csa_tree_add_48_2_groupi_n_1196 & ~n_179) | (csa_tree_add_48_2_groupi_n_1305
    & n_179));
 assign csa_tree_add_48_2_groupi_n_1348 = ~(csa_tree_add_48_2_groupi_n_1297 ^ csa_tree_add_48_2_groupi_n_979);
 assign csa_tree_add_48_2_groupi_n_1359 = ~(csa_tree_add_48_2_groupi_n_1329 | csa_tree_add_48_2_groupi_n_1330);
 assign csa_tree_add_48_2_groupi_n_1347 = ~(csa_tree_add_48_2_groupi_n_1326 & ~(csa_tree_add_48_2_groupi_n_1304
    & csa_tree_add_48_2_groupi_n_1272));
 assign csa_tree_add_48_2_groupi_n_1341 = ~((csa_tree_add_48_2_groupi_n_1195 & ~csa_tree_add_48_2_groupi_n_1308)
    | (csa_tree_add_48_2_groupi_n_1303 & csa_tree_add_48_2_groupi_n_1308));
 assign csa_tree_add_48_2_groupi_n_1346 = ~(csa_tree_add_48_2_groupi_n_1331 | csa_tree_add_48_2_groupi_n_1332);
 assign csa_tree_add_48_2_groupi_n_1340 = ~((csa_tree_add_48_2_groupi_n_1300 & ~csa_tree_add_48_2_groupi_n_1312)
    | (csa_tree_add_48_2_groupi_n_1192 & csa_tree_add_48_2_groupi_n_1312));
 assign csa_tree_add_48_2_groupi_n_1345 = ~(csa_tree_add_48_2_groupi_n_1317 & csa_tree_add_48_2_groupi_n_1155);
 assign csa_tree_add_48_2_groupi_n_1339 = ~(csa_tree_add_48_2_groupi_n_1325 & csa_tree_add_48_2_groupi_n_1136);
 assign csa_tree_add_48_2_groupi_n_1338 = ~(csa_tree_add_48_2_groupi_n_1156 & (csa_tree_add_48_2_groupi_n_1153
    | csa_tree_add_48_2_groupi_n_1157));
 assign csa_tree_add_48_2_groupi_n_1336 = (csa_tree_add_48_2_groupi_n_1167 & csa_tree_add_48_2_groupi_n_749);
 assign csa_tree_add_48_2_groupi_n_1337 = (csa_tree_add_48_2_groupi_n_1167 ^ csa_tree_add_48_2_groupi_n_749);
 assign csa_tree_add_48_2_groupi_n_1335 = ~(n_178 & csa_tree_add_48_2_groupi_n_1128);
 assign csa_tree_add_48_2_groupi_n_1334 = ~(csa_tree_add_48_2_groupi_n_1314 & csa_tree_add_48_2_groupi_n_1315);
 assign csa_tree_add_48_2_groupi_n_1333 = ~(csa_tree_add_48_2_groupi_n_1314 | csa_tree_add_48_2_groupi_n_1315);
 assign csa_tree_add_48_2_groupi_n_1332 = ~(n_178 | n_182);
 assign csa_tree_add_48_2_groupi_n_1331 = ~(csa_tree_add_48_2_groupi_n_1299 | csa_tree_add_48_2_groupi_n_1128);
 assign csa_tree_add_48_2_groupi_n_1330 = ~(csa_tree_add_48_2_groupi_n_1277 | csa_tree_add_48_2_groupi_n_1314);
 assign csa_tree_add_48_2_groupi_n_1329 = ~(csa_tree_add_48_2_groupi_n_1278 | csa_tree_add_48_2_groupi_n_1190);
 assign csa_tree_add_48_2_groupi_n_1328 = ~(csa_tree_add_48_2_groupi_n_1312 | csa_tree_add_48_2_groupi_n_1300);
 assign csa_tree_add_48_2_groupi_n_1325 = ~(csa_tree_add_48_2_groupi_n_1138 & ~csa_tree_add_48_2_groupi_n_135);
 assign csa_tree_add_48_2_groupi_n_1324 = ~(csa_tree_add_48_2_groupi_n_1276 | csa_tree_add_48_2_groupi_n_1313);
 assign csa_tree_add_48_2_groupi_n_1323 = ~(csa_tree_add_48_2_groupi_n_35 | n_179);
 assign csa_tree_add_48_2_groupi_n_1322 = ~(csa_tree_add_48_2_groupi_n_35 & n_179);
 assign csa_tree_add_48_2_groupi_n_1321 = ~(csa_tree_add_48_2_groupi_n_1189 & csa_tree_add_48_2_groupi_n_1268);
 assign csa_tree_add_48_2_groupi_n_1320 = ~(csa_tree_add_48_2_groupi_n_1299 & n_182);
 assign csa_tree_add_48_2_groupi_n_1319 = ~(csa_tree_add_48_2_groupi_n_1312 & csa_tree_add_48_2_groupi_n_1300);
 assign csa_tree_add_48_2_groupi_n_1318 = ~(csa_tree_add_48_2_groupi_n_1276 & csa_tree_add_48_2_groupi_n_1313);
 assign csa_tree_add_48_2_groupi_n_1317 = ~(csa_tree_add_48_2_groupi_n_1275 & csa_tree_add_48_2_groupi_n_1160);
 assign csa_tree_add_48_2_groupi_n_1326 = (csa_tree_add_48_2_groupi_n_1304 | csa_tree_add_48_2_groupi_n_1272);
 assign csa_tree_add_48_2_groupi_n_1314 = ~csa_tree_add_48_2_groupi_n_1190;
 assign csa_tree_add_48_2_groupi_n_1309 = ~csa_tree_add_48_2_groupi_n_1194;
 assign csa_tree_add_48_2_groupi_n_1305 = ~csa_tree_add_48_2_groupi_n_1196;
 assign csa_tree_add_48_2_groupi_n_1303 = ~csa_tree_add_48_2_groupi_n_1195;
 assign csa_tree_add_48_2_groupi_n_1301 = ~csa_tree_add_48_2_groupi_n_1302;
 assign csa_tree_add_48_2_groupi_n_1300 = ~csa_tree_add_48_2_groupi_n_1192;
 assign csa_tree_add_48_2_groupi_n_1299 = ~n_178;
 assign csa_tree_add_48_2_groupi_n_1297 = ((csa_tree_add_48_2_groupi_n_909 & csa_tree_add_48_2_groupi_n_954)
    | ((csa_tree_add_48_2_groupi_n_954 & csa_tree_add_48_2_groupi_n_1058) | (csa_tree_add_48_2_groupi_n_1058
    & csa_tree_add_48_2_groupi_n_909)));
 assign csa_tree_add_48_2_groupi_n_1298 = (csa_tree_add_48_2_groupi_n_954 ^ (csa_tree_add_48_2_groupi_n_1058
    ^ csa_tree_add_48_2_groupi_n_909));
 assign csa_tree_add_48_2_groupi_n_1315 = ((csa_tree_add_48_2_groupi_n_907 & csa_tree_add_48_2_groupi_n_1039)
    | ((csa_tree_add_48_2_groupi_n_1039 & csa_tree_add_48_2_groupi_n_1056) | (csa_tree_add_48_2_groupi_n_1056
    & csa_tree_add_48_2_groupi_n_907)));
 assign csa_tree_add_48_2_groupi_n_1316 = (csa_tree_add_48_2_groupi_n_1039 ^ (csa_tree_add_48_2_groupi_n_1056
    ^ csa_tree_add_48_2_groupi_n_907));
 assign csa_tree_add_48_2_groupi_n_1295 = ((csa_tree_add_48_2_groupi_n_882 & csa_tree_add_48_2_groupi_n_952)
    | ((csa_tree_add_48_2_groupi_n_952 & csa_tree_add_48_2_groupi_n_1035) | (csa_tree_add_48_2_groupi_n_1035
    & csa_tree_add_48_2_groupi_n_882)));
 assign csa_tree_add_48_2_groupi_n_1296 = (csa_tree_add_48_2_groupi_n_952 ^ (csa_tree_add_48_2_groupi_n_1035
    ^ csa_tree_add_48_2_groupi_n_882));
 assign csa_tree_add_48_2_groupi_n_1312 = ((csa_tree_add_48_2_groupi_n_966 & csa_tree_add_48_2_groupi_n_1055)
    | ((csa_tree_add_48_2_groupi_n_1055 & csa_tree_add_48_2_groupi_n_960) | (csa_tree_add_48_2_groupi_n_960
    & csa_tree_add_48_2_groupi_n_966)));
 assign csa_tree_add_48_2_groupi_n_1313 = (csa_tree_add_48_2_groupi_n_1055 ^ (csa_tree_add_48_2_groupi_n_960
    ^ csa_tree_add_48_2_groupi_n_966));
 assign csa_tree_add_48_2_groupi_n_1310 = ((csa_tree_add_48_2_groupi_n_1040 & csa_tree_add_48_2_groupi_n_1057)
    | ((csa_tree_add_48_2_groupi_n_1057 & csa_tree_add_48_2_groupi_n_1054) | (csa_tree_add_48_2_groupi_n_1054
    & csa_tree_add_48_2_groupi_n_1040)));
 assign csa_tree_add_48_2_groupi_n_1311 = (csa_tree_add_48_2_groupi_n_1057 ^ (csa_tree_add_48_2_groupi_n_1054
    ^ csa_tree_add_48_2_groupi_n_1040));
 assign csa_tree_add_48_2_groupi_n_1307 = ((csa_tree_add_48_2_groupi_n_1042 & csa_tree_add_48_2_groupi_n_963)
    | ((csa_tree_add_48_2_groupi_n_963 & csa_tree_add_48_2_groupi_n_1053) | (csa_tree_add_48_2_groupi_n_1053
    & csa_tree_add_48_2_groupi_n_1042)));
 assign csa_tree_add_48_2_groupi_n_1308 = (csa_tree_add_48_2_groupi_n_963 ^ (csa_tree_add_48_2_groupi_n_1053
    ^ csa_tree_add_48_2_groupi_n_1042));
 assign csa_tree_add_48_2_groupi_n_1294 = ((csa_tree_add_48_2_groupi_n_900 & csa_tree_add_48_2_groupi_n_1033)
    | ((csa_tree_add_48_2_groupi_n_1033 & csa_tree_add_48_2_groupi_n_864) | (csa_tree_add_48_2_groupi_n_864
    & csa_tree_add_48_2_groupi_n_900)));
 assign csa_tree_add_48_2_groupi_n_1304 = (csa_tree_add_48_2_groupi_n_1033 ^ (csa_tree_add_48_2_groupi_n_864
    ^ csa_tree_add_48_2_groupi_n_900));
 assign csa_tree_add_48_2_groupi_n_1292 = ((csa_tree_add_48_2_groupi_n_901 & csa_tree_add_48_2_groupi_n_1029)
    | ((csa_tree_add_48_2_groupi_n_1029 & csa_tree_add_48_2_groupi_n_868) | (csa_tree_add_48_2_groupi_n_868
    & csa_tree_add_48_2_groupi_n_901)));
 assign csa_tree_add_48_2_groupi_n_1293 = (csa_tree_add_48_2_groupi_n_1029 ^ (csa_tree_add_48_2_groupi_n_868
    ^ csa_tree_add_48_2_groupi_n_901));
 assign csa_tree_add_48_2_groupi_n_1290 = ((csa_tree_add_48_2_groupi_n_888 & csa_tree_add_48_2_groupi_n_1027)
    | ((csa_tree_add_48_2_groupi_n_1027 & csa_tree_add_48_2_groupi_n_869) | (csa_tree_add_48_2_groupi_n_869
    & csa_tree_add_48_2_groupi_n_888)));
 assign csa_tree_add_48_2_groupi_n_1291 = (csa_tree_add_48_2_groupi_n_1027 ^ (csa_tree_add_48_2_groupi_n_869
    ^ csa_tree_add_48_2_groupi_n_888));
 assign csa_tree_add_48_2_groupi_n_1289 = ((csa_tree_add_48_2_groupi_n_967 & csa_tree_add_48_2_groupi_n_1060)
    | ((csa_tree_add_48_2_groupi_n_1060 & csa_tree_add_48_2_groupi_n_956) | (csa_tree_add_48_2_groupi_n_956
    & csa_tree_add_48_2_groupi_n_967)));
 assign csa_tree_add_48_2_groupi_n_1302 = (csa_tree_add_48_2_groupi_n_1060 ^ (csa_tree_add_48_2_groupi_n_956
    ^ csa_tree_add_48_2_groupi_n_967));
 assign csa_tree_add_48_2_groupi_n_1287 = ((csa_tree_add_48_2_groupi_n_908 & csa_tree_add_48_2_groupi_n_1052)
    | ((csa_tree_add_48_2_groupi_n_1052 & csa_tree_add_48_2_groupi_n_1037) | (csa_tree_add_48_2_groupi_n_1037
    & csa_tree_add_48_2_groupi_n_908)));
 assign csa_tree_add_48_2_groupi_n_1288 = (csa_tree_add_48_2_groupi_n_1052 ^ (csa_tree_add_48_2_groupi_n_1037
    ^ csa_tree_add_48_2_groupi_n_908));
 assign csa_tree_add_48_2_groupi_n_1285 = ((csa_tree_add_48_2_groupi_n_903 & csa_tree_add_48_2_groupi_n_1036)
    | ((csa_tree_add_48_2_groupi_n_1036 & csa_tree_add_48_2_groupi_n_866) | (csa_tree_add_48_2_groupi_n_866
    & csa_tree_add_48_2_groupi_n_903)));
 assign csa_tree_add_48_2_groupi_n_1286 = (csa_tree_add_48_2_groupi_n_1036 ^ (csa_tree_add_48_2_groupi_n_866
    ^ csa_tree_add_48_2_groupi_n_903));
 assign csa_tree_add_48_2_groupi_n_1284 = ~((csa_tree_add_48_2_groupi_n_1070 & ~csa_tree_add_48_2_groupi_n_1115)
    | (csa_tree_add_48_2_groupi_n_132 & csa_tree_add_48_2_groupi_n_1115));
 assign csa_tree_add_48_2_groupi_n_1283 = ~((csa_tree_add_48_2_groupi_n_1046 & ~csa_tree_add_48_2_groupi_n_1183)
    | (csa_tree_add_48_2_groupi_n_1127 & csa_tree_add_48_2_groupi_n_1183));
 assign csa_tree_add_48_2_groupi_n_1282 = ~((csa_tree_add_48_2_groupi_n_1181 & ~csa_tree_add_48_2_groupi_n_22)
    | (csa_tree_add_48_2_groupi_n_1182 & csa_tree_add_48_2_groupi_n_22));
 assign csa_tree_add_48_2_groupi_n_1278 = ~csa_tree_add_48_2_groupi_n_1277;
 assign csa_tree_add_48_2_groupi_n_1267 = ((csa_tree_add_48_2_groupi_n_902 & csa_tree_add_48_2_groupi_n_308)
    | ((csa_tree_add_48_2_groupi_n_308 & csa_tree_add_48_2_groupi_n_949) | (csa_tree_add_48_2_groupi_n_949
    & csa_tree_add_48_2_groupi_n_902)));
 assign csa_tree_add_48_2_groupi_n_1281 = (csa_tree_add_48_2_groupi_n_308 ^ (csa_tree_add_48_2_groupi_n_949
    ^ csa_tree_add_48_2_groupi_n_902));
 assign csa_tree_add_48_2_groupi_n_1265 = ((csa_tree_add_48_2_groupi_n_880 & csa_tree_add_48_2_groupi_n_312)
    | ((csa_tree_add_48_2_groupi_n_312 & csa_tree_add_48_2_groupi_n_856) | (csa_tree_add_48_2_groupi_n_856
    & csa_tree_add_48_2_groupi_n_880)));
 assign csa_tree_add_48_2_groupi_n_1266 = (csa_tree_add_48_2_groupi_n_312 ^ (csa_tree_add_48_2_groupi_n_856
    ^ csa_tree_add_48_2_groupi_n_880));
 assign csa_tree_add_48_2_groupi_n_1277 = ((csa_tree_add_48_2_groupi_n_887 & csa_tree_add_48_2_groupi_n_964)
    | ((csa_tree_add_48_2_groupi_n_964 & csa_tree_add_48_2_groupi_n_948) | (csa_tree_add_48_2_groupi_n_948
    & csa_tree_add_48_2_groupi_n_887)));
 assign csa_tree_add_48_2_groupi_n_1280 = (csa_tree_add_48_2_groupi_n_964 ^ (csa_tree_add_48_2_groupi_n_948
    ^ csa_tree_add_48_2_groupi_n_887));
 assign csa_tree_add_48_2_groupi_n_1263 = ((csa_tree_add_48_2_groupi_n_928 & csa_tree_add_48_2_groupi_n_1034)
    | ((csa_tree_add_48_2_groupi_n_1034 & csa_tree_add_48_2_groupi_n_925) | (csa_tree_add_48_2_groupi_n_925
    & csa_tree_add_48_2_groupi_n_928)));
 assign csa_tree_add_48_2_groupi_n_1264 = (csa_tree_add_48_2_groupi_n_1034 ^ (csa_tree_add_48_2_groupi_n_925
    ^ csa_tree_add_48_2_groupi_n_928));
 assign csa_tree_add_48_2_groupi_n_1261 = ((csa_tree_add_48_2_groupi_n_997 & csa_tree_add_48_2_groupi_n_1022)
    | ((csa_tree_add_48_2_groupi_n_1022 & csa_tree_add_48_2_groupi_n_921) | (csa_tree_add_48_2_groupi_n_921
    & csa_tree_add_48_2_groupi_n_997)));
 assign csa_tree_add_48_2_groupi_n_1262 = (csa_tree_add_48_2_groupi_n_1022 ^ (csa_tree_add_48_2_groupi_n_921
    ^ csa_tree_add_48_2_groupi_n_997));
 assign csa_tree_add_48_2_groupi_n_1259 = ((csa_tree_add_48_2_groupi_n_890 & csa_tree_add_48_2_groupi_n_324)
    | ((csa_tree_add_48_2_groupi_n_324 & csa_tree_add_48_2_groupi_n_863) | (csa_tree_add_48_2_groupi_n_863
    & csa_tree_add_48_2_groupi_n_890)));
 assign csa_tree_add_48_2_groupi_n_1260 = (csa_tree_add_48_2_groupi_n_324 ^ (csa_tree_add_48_2_groupi_n_863
    ^ csa_tree_add_48_2_groupi_n_890));
 assign csa_tree_add_48_2_groupi_n_1275 = ((csa_tree_add_48_2_groupi_n_881 & csa_tree_add_48_2_groupi_n_962)
    | ((csa_tree_add_48_2_groupi_n_962 & csa_tree_add_48_2_groupi_n_961) | (csa_tree_add_48_2_groupi_n_961
    & csa_tree_add_48_2_groupi_n_881)));
 assign csa_tree_add_48_2_groupi_n_1276 = (csa_tree_add_48_2_groupi_n_962 ^ (csa_tree_add_48_2_groupi_n_961
    ^ csa_tree_add_48_2_groupi_n_881));
 assign csa_tree_add_48_2_groupi_n_1257 = ((csa_tree_add_48_2_groupi_n_999 & csa_tree_add_48_2_groupi_n_1059)
    | ((csa_tree_add_48_2_groupi_n_1059 & csa_tree_add_48_2_groupi_n_996) | (csa_tree_add_48_2_groupi_n_996
    & csa_tree_add_48_2_groupi_n_999)));
 assign csa_tree_add_48_2_groupi_n_1258 = (csa_tree_add_48_2_groupi_n_1059 ^ (csa_tree_add_48_2_groupi_n_996
    ^ csa_tree_add_48_2_groupi_n_999));
 assign csa_tree_add_48_2_groupi_n_1255 = ((csa_tree_add_48_2_groupi_n_879 & csa_tree_add_48_2_groupi_n_714)
    | ((csa_tree_add_48_2_groupi_n_714 & csa_tree_add_48_2_groupi_n_950) | (csa_tree_add_48_2_groupi_n_950
    & csa_tree_add_48_2_groupi_n_879)));
 assign csa_tree_add_48_2_groupi_n_1256 = (csa_tree_add_48_2_groupi_n_714 ^ (csa_tree_add_48_2_groupi_n_950
    ^ csa_tree_add_48_2_groupi_n_879));
 assign csa_tree_add_48_2_groupi_n_1253 = ((csa_tree_add_48_2_groupi_n_924 & csa_tree_add_48_2_groupi_n_1030)
    | ((csa_tree_add_48_2_groupi_n_1030 & csa_tree_add_48_2_groupi_n_931) | (csa_tree_add_48_2_groupi_n_931
    & csa_tree_add_48_2_groupi_n_924)));
 assign csa_tree_add_48_2_groupi_n_1254 = (csa_tree_add_48_2_groupi_n_1030 ^ (csa_tree_add_48_2_groupi_n_931
    ^ csa_tree_add_48_2_groupi_n_924));
 assign csa_tree_add_48_2_groupi_n_1251 = ((csa_tree_add_48_2_groupi_n_926 & csa_tree_add_48_2_groupi_n_1032)
    | ((csa_tree_add_48_2_groupi_n_1032 & csa_tree_add_48_2_groupi_n_913) | (csa_tree_add_48_2_groupi_n_913
    & csa_tree_add_48_2_groupi_n_926)));
 assign csa_tree_add_48_2_groupi_n_1252 = (csa_tree_add_48_2_groupi_n_1032 ^ (csa_tree_add_48_2_groupi_n_913
    ^ csa_tree_add_48_2_groupi_n_926));
 assign csa_tree_add_48_2_groupi_n_1249 = ((csa_tree_add_48_2_groupi_n_891 & csa_tree_add_48_2_groupi_n_323)
    | ((csa_tree_add_48_2_groupi_n_323 & csa_tree_add_48_2_groupi_n_874) | (csa_tree_add_48_2_groupi_n_874
    & csa_tree_add_48_2_groupi_n_891)));
 assign csa_tree_add_48_2_groupi_n_1250 = (csa_tree_add_48_2_groupi_n_323 ^ (csa_tree_add_48_2_groupi_n_874
    ^ csa_tree_add_48_2_groupi_n_891));
 assign csa_tree_add_48_2_groupi_n_1247 = ((csa_tree_add_48_2_groupi_n_893 & csa_tree_add_48_2_groupi_n_314)
    | ((csa_tree_add_48_2_groupi_n_314 & csa_tree_add_48_2_groupi_n_870) | (csa_tree_add_48_2_groupi_n_870
    & csa_tree_add_48_2_groupi_n_893)));
 assign csa_tree_add_48_2_groupi_n_1248 = (csa_tree_add_48_2_groupi_n_314 ^ (csa_tree_add_48_2_groupi_n_870
    ^ csa_tree_add_48_2_groupi_n_893));
 assign csa_tree_add_48_2_groupi_n_1245 = ((csa_tree_add_48_2_groupi_n_886 & csa_tree_add_48_2_groupi_n_1061)
    | ((csa_tree_add_48_2_groupi_n_1061 & csa_tree_add_48_2_groupi_n_1043) | (csa_tree_add_48_2_groupi_n_1043
    & csa_tree_add_48_2_groupi_n_886)));
 assign csa_tree_add_48_2_groupi_n_1246 = (csa_tree_add_48_2_groupi_n_1061 ^ (csa_tree_add_48_2_groupi_n_1043
    ^ csa_tree_add_48_2_groupi_n_886));
 assign csa_tree_add_48_2_groupi_n_1243 = ((csa_tree_add_48_2_groupi_n_885 & csa_tree_add_48_2_groupi_n_317)
    | ((csa_tree_add_48_2_groupi_n_317 & csa_tree_add_48_2_groupi_n_867) | (csa_tree_add_48_2_groupi_n_867
    & csa_tree_add_48_2_groupi_n_885)));
 assign csa_tree_add_48_2_groupi_n_1244 = (csa_tree_add_48_2_groupi_n_317 ^ (csa_tree_add_48_2_groupi_n_867
    ^ csa_tree_add_48_2_groupi_n_885));
 assign csa_tree_add_48_2_groupi_n_1242 = ((csa_tree_add_48_2_groupi_n_968 & csa_tree_add_48_2_groupi_n_325)
    | ((csa_tree_add_48_2_groupi_n_325 & csa_tree_add_48_2_groupi_n_24) | (csa_tree_add_48_2_groupi_n_24
    & csa_tree_add_48_2_groupi_n_968)));
 assign csa_tree_add_48_2_groupi_n_1274 = (csa_tree_add_48_2_groupi_n_325 ^ (csa_tree_add_48_2_groupi_n_24
    ^ csa_tree_add_48_2_groupi_n_968));
 assign csa_tree_add_48_2_groupi_n_1240 = ((csa_tree_add_48_2_groupi_n_894 & csa_tree_add_48_2_groupi_n_320)
    | ((csa_tree_add_48_2_groupi_n_320 & csa_tree_add_48_2_groupi_n_857) | (csa_tree_add_48_2_groupi_n_857
    & csa_tree_add_48_2_groupi_n_894)));
 assign csa_tree_add_48_2_groupi_n_1241 = (csa_tree_add_48_2_groupi_n_320 ^ (csa_tree_add_48_2_groupi_n_857
    ^ csa_tree_add_48_2_groupi_n_894));
 assign csa_tree_add_48_2_groupi_n_1238 = ((csa_tree_add_48_2_groupi_n_910 & csa_tree_add_48_2_groupi_n_326)
    | ((csa_tree_add_48_2_groupi_n_326 & csa_tree_add_48_2_groupi_n_861) | (csa_tree_add_48_2_groupi_n_861
    & csa_tree_add_48_2_groupi_n_910)));
 assign csa_tree_add_48_2_groupi_n_1239 = (csa_tree_add_48_2_groupi_n_326 ^ (csa_tree_add_48_2_groupi_n_861
    ^ csa_tree_add_48_2_groupi_n_910));
 assign csa_tree_add_48_2_groupi_n_1236 = ((csa_tree_add_48_2_groupi_n_969 & csa_tree_add_48_2_groupi_n_951)
    | ((csa_tree_add_48_2_groupi_n_951 & csa_tree_add_48_2_groupi_n_957) | (csa_tree_add_48_2_groupi_n_957
    & csa_tree_add_48_2_groupi_n_969)));
 assign csa_tree_add_48_2_groupi_n_1237 = (csa_tree_add_48_2_groupi_n_951 ^ (csa_tree_add_48_2_groupi_n_957
    ^ csa_tree_add_48_2_groupi_n_969));
 assign csa_tree_add_48_2_groupi_n_1234 = ((csa_tree_add_48_2_groupi_n_922 & csa_tree_add_48_2_groupi_n_1023)
    | ((csa_tree_add_48_2_groupi_n_1023 & csa_tree_add_48_2_groupi_n_933) | (csa_tree_add_48_2_groupi_n_933
    & csa_tree_add_48_2_groupi_n_922)));
 assign csa_tree_add_48_2_groupi_n_1235 = (csa_tree_add_48_2_groupi_n_1023 ^ (csa_tree_add_48_2_groupi_n_933
    ^ csa_tree_add_48_2_groupi_n_922));
 assign csa_tree_add_48_2_groupi_n_1233 = ((csa_tree_add_48_2_groupi_n_977 & csa_tree_add_48_2_groupi_n_26)
    | ((csa_tree_add_48_2_groupi_n_26 & csa_tree_add_48_2_groupi_n_958) | (csa_tree_add_48_2_groupi_n_958
    & csa_tree_add_48_2_groupi_n_977)));
 assign csa_tree_add_48_2_groupi_n_1273 = (csa_tree_add_48_2_groupi_n_26 ^ (csa_tree_add_48_2_groupi_n_958
    ^ csa_tree_add_48_2_groupi_n_977));
 assign csa_tree_add_48_2_groupi_n_1231 = ((csa_tree_add_48_2_groupi_n_883 & csa_tree_add_48_2_groupi_n_319)
    | ((csa_tree_add_48_2_groupi_n_319 & csa_tree_add_48_2_groupi_n_873) | (csa_tree_add_48_2_groupi_n_873
    & csa_tree_add_48_2_groupi_n_883)));
 assign csa_tree_add_48_2_groupi_n_1232 = (csa_tree_add_48_2_groupi_n_319 ^ (csa_tree_add_48_2_groupi_n_873
    ^ csa_tree_add_48_2_groupi_n_883));
 assign csa_tree_add_48_2_groupi_n_1229 = ((csa_tree_add_48_2_groupi_n_932 & csa_tree_add_48_2_groupi_n_1026)
    | ((csa_tree_add_48_2_groupi_n_1026 & csa_tree_add_48_2_groupi_n_935) | (csa_tree_add_48_2_groupi_n_935
    & csa_tree_add_48_2_groupi_n_932)));
 assign csa_tree_add_48_2_groupi_n_1230 = (csa_tree_add_48_2_groupi_n_1026 ^ (csa_tree_add_48_2_groupi_n_935
    ^ csa_tree_add_48_2_groupi_n_932));
 assign csa_tree_add_48_2_groupi_n_1272 = ((csa_tree_add_48_2_groupi_n_905 & csa_tree_add_48_2_groupi_n_328)
    | ((csa_tree_add_48_2_groupi_n_328 & csa_tree_add_48_2_groupi_n_1028) | (csa_tree_add_48_2_groupi_n_1028
    & csa_tree_add_48_2_groupi_n_905)));
 assign csa_tree_add_48_2_groupi_n_1228 = (csa_tree_add_48_2_groupi_n_328 ^ (csa_tree_add_48_2_groupi_n_1028
    ^ csa_tree_add_48_2_groupi_n_905));
 assign csa_tree_add_48_2_groupi_n_1226 = ((csa_tree_add_48_2_groupi_n_889 & csa_tree_add_48_2_groupi_n_310)
    | ((csa_tree_add_48_2_groupi_n_310 & csa_tree_add_48_2_groupi_n_860) | (csa_tree_add_48_2_groupi_n_860
    & csa_tree_add_48_2_groupi_n_889)));
 assign csa_tree_add_48_2_groupi_n_1227 = (csa_tree_add_48_2_groupi_n_310 ^ (csa_tree_add_48_2_groupi_n_860
    ^ csa_tree_add_48_2_groupi_n_889));
 assign csa_tree_add_48_2_groupi_n_1224 = ((csa_tree_add_48_2_groupi_n_936 & csa_tree_add_48_2_groupi_n_1021)
    | ((csa_tree_add_48_2_groupi_n_1021 & csa_tree_add_48_2_groupi_n_929) | (csa_tree_add_48_2_groupi_n_929
    & csa_tree_add_48_2_groupi_n_936)));
 assign csa_tree_add_48_2_groupi_n_1225 = (csa_tree_add_48_2_groupi_n_1021 ^ (csa_tree_add_48_2_groupi_n_929
    ^ csa_tree_add_48_2_groupi_n_936));
 assign csa_tree_add_48_2_groupi_n_1223 = ((csa_tree_add_48_2_groupi_n_898 & csa_tree_add_48_2_groupi_n_959)
    | ((csa_tree_add_48_2_groupi_n_959 & csa_tree_add_48_2_groupi_n_878) | (csa_tree_add_48_2_groupi_n_878
    & csa_tree_add_48_2_groupi_n_898)));
 assign csa_tree_add_48_2_groupi_n_1271 = (csa_tree_add_48_2_groupi_n_959 ^ (csa_tree_add_48_2_groupi_n_878
    ^ csa_tree_add_48_2_groupi_n_898));
 assign csa_tree_add_48_2_groupi_n_1221 = ((csa_tree_add_48_2_groupi_n_906 & csa_tree_add_48_2_groupi_n_1025)
    | ((csa_tree_add_48_2_groupi_n_1025 & csa_tree_add_48_2_groupi_n_875) | (csa_tree_add_48_2_groupi_n_875
    & csa_tree_add_48_2_groupi_n_906)));
 assign csa_tree_add_48_2_groupi_n_1222 = (csa_tree_add_48_2_groupi_n_1025 ^ (csa_tree_add_48_2_groupi_n_875
    ^ csa_tree_add_48_2_groupi_n_906));
 assign csa_tree_add_48_2_groupi_n_1219 = ((csa_tree_add_48_2_groupi_n_971 & csa_tree_add_48_2_groupi_n_872)
    | ((csa_tree_add_48_2_groupi_n_872 & csa_tree_add_48_2_groupi_n_309) | (csa_tree_add_48_2_groupi_n_309
    & csa_tree_add_48_2_groupi_n_971)));
 assign csa_tree_add_48_2_groupi_n_1220 = (csa_tree_add_48_2_groupi_n_872 ^ (csa_tree_add_48_2_groupi_n_309
    ^ csa_tree_add_48_2_groupi_n_971));
 assign csa_tree_add_48_2_groupi_n_1217 = ((csa_tree_add_48_2_groupi_n_897 & csa_tree_add_48_2_groupi_n_321)
    | ((csa_tree_add_48_2_groupi_n_321 & csa_tree_add_48_2_groupi_n_859) | (csa_tree_add_48_2_groupi_n_859
    & csa_tree_add_48_2_groupi_n_897)));
 assign csa_tree_add_48_2_groupi_n_1218 = (csa_tree_add_48_2_groupi_n_321 ^ (csa_tree_add_48_2_groupi_n_859
    ^ csa_tree_add_48_2_groupi_n_897));
 assign csa_tree_add_48_2_groupi_n_1215 = ((csa_tree_add_48_2_groupi_n_904 & csa_tree_add_48_2_groupi_n_953)
    | ((csa_tree_add_48_2_groupi_n_953 & csa_tree_add_48_2_groupi_n_865) | (csa_tree_add_48_2_groupi_n_865
    & csa_tree_add_48_2_groupi_n_904)));
 assign csa_tree_add_48_2_groupi_n_1216 = (csa_tree_add_48_2_groupi_n_953 ^ (csa_tree_add_48_2_groupi_n_865
    ^ csa_tree_add_48_2_groupi_n_904));
 assign csa_tree_add_48_2_groupi_n_1213 = ((csa_tree_add_48_2_groupi_n_911 & csa_tree_add_48_2_groupi_n_871)
    | ((csa_tree_add_48_2_groupi_n_871 & csa_tree_add_48_2_groupi_n_955) | (csa_tree_add_48_2_groupi_n_955
    & csa_tree_add_48_2_groupi_n_911)));
 assign csa_tree_add_48_2_groupi_n_1214 = (csa_tree_add_48_2_groupi_n_871 ^ (csa_tree_add_48_2_groupi_n_955
    ^ csa_tree_add_48_2_groupi_n_911));
 assign csa_tree_add_48_2_groupi_n_1211 = ((csa_tree_add_48_2_groupi_n_934 & csa_tree_add_48_2_groupi_n_1024)
    | ((csa_tree_add_48_2_groupi_n_1024 & csa_tree_add_48_2_groupi_n_923) | (csa_tree_add_48_2_groupi_n_923
    & csa_tree_add_48_2_groupi_n_934)));
 assign csa_tree_add_48_2_groupi_n_1212 = (csa_tree_add_48_2_groupi_n_1024 ^ (csa_tree_add_48_2_groupi_n_923
    ^ csa_tree_add_48_2_groupi_n_934));
 assign csa_tree_add_48_2_groupi_n_1209 = ((csa_tree_add_48_2_groupi_n_892 & csa_tree_add_48_2_groupi_n_318)
    | ((csa_tree_add_48_2_groupi_n_318 & csa_tree_add_48_2_groupi_n_858) | (csa_tree_add_48_2_groupi_n_858
    & csa_tree_add_48_2_groupi_n_892)));
 assign csa_tree_add_48_2_groupi_n_1210 = (csa_tree_add_48_2_groupi_n_318 ^ (csa_tree_add_48_2_groupi_n_858
    ^ csa_tree_add_48_2_groupi_n_892));
 assign csa_tree_add_48_2_groupi_n_1207 = ((csa_tree_add_48_2_groupi_n_930 & csa_tree_add_48_2_groupi_n_1031)
    | ((csa_tree_add_48_2_groupi_n_1031 & csa_tree_add_48_2_groupi_n_927) | (csa_tree_add_48_2_groupi_n_927
    & csa_tree_add_48_2_groupi_n_930)));
 assign csa_tree_add_48_2_groupi_n_1208 = (csa_tree_add_48_2_groupi_n_1031 ^ (csa_tree_add_48_2_groupi_n_927
    ^ csa_tree_add_48_2_groupi_n_930));
 assign csa_tree_add_48_2_groupi_n_1206 = ~(csa_tree_add_48_2_groupi_n_1184 & ~csa_tree_add_48_2_groupi_n_1046);
 assign csa_tree_add_48_2_groupi_n_1205 = ~(csa_tree_add_48_2_groupi_n_23 | csa_tree_add_48_2_groupi_n_1135);
 assign csa_tree_add_48_2_groupi_n_1204 = ~(n_180 & csa_tree_add_48_2_groupi_n_1124);
 assign csa_tree_add_48_2_groupi_n_1203 = ~(csa_tree_add_48_2_groupi_n_1115 | csa_tree_add_48_2_groupi_n_1070);
 assign csa_tree_add_48_2_groupi_n_1202 = ~(csa_tree_add_48_2_groupi_n_1131 & csa_tree_add_48_2_groupi_n_1182);
 assign csa_tree_add_48_2_groupi_n_1201 = ~(csa_tree_add_48_2_groupi_n_23 & csa_tree_add_48_2_groupi_n_1135);
 assign csa_tree_add_48_2_groupi_n_1200 = ~(csa_tree_add_48_2_groupi_n_1184 | csa_tree_add_48_2_groupi_n_1127);
 assign csa_tree_add_48_2_groupi_n_1199 = ~(n_180 | csa_tree_add_48_2_groupi_n_1124);
 assign csa_tree_add_48_2_groupi_n_1270 = ~(csa_tree_add_48_2_groupi_n_1158 | csa_tree_add_48_2_groupi_n_1159);
 assign csa_tree_add_48_2_groupi_n_135 = ~(csa_tree_add_48_2_groupi_n_1110 | (csa_tree_add_48_2_groupi_n_1094
    & csa_tree_add_48_2_groupi_n_1050));
 assign csa_tree_add_48_2_groupi_n_1198 = ~(csa_tree_add_48_2_groupi_n_1151 & csa_tree_add_48_2_groupi_n_1109);
 assign csa_tree_add_48_2_groupi_n_1268 = ~(csa_tree_add_48_2_groupi_n_1111 & (csa_tree_add_48_2_groupi_n_1095
    | csa_tree_add_48_2_groupi_n_941));
 assign csa_tree_add_48_2_groupi_n_1197 = ~(csa_tree_add_48_2_groupi_n_1112 ^ csa_tree_add_48_2_groupi_n_938);
 assign csa_tree_add_48_2_groupi_n_1196 = ~(csa_tree_add_48_2_groupi_n_1147 | csa_tree_add_48_2_groupi_n_44);
 assign csa_tree_add_48_2_groupi_n_1195 = ~(csa_tree_add_48_2_groupi_n_1146 | csa_tree_add_48_2_groupi_n_43);
 assign csa_tree_add_48_2_groupi_n_1194 = ~(csa_tree_add_48_2_groupi_n_1149 | csa_tree_add_48_2_groupi_n_1102);
 assign csa_tree_add_48_2_groupi_n_1193 = ~(csa_tree_add_48_2_groupi_n_1145 | csa_tree_add_48_2_groupi_n_1100);
 assign csa_tree_add_48_2_groupi_n_1192 = ~(csa_tree_add_48_2_groupi_n_1148 | csa_tree_add_48_2_groupi_n_1107);
 assign csa_tree_add_48_2_groupi_n_1186 = ~(csa_tree_add_48_2_groupi_n_1106 & (csa_tree_add_48_2_groupi_n_1105
    | csa_tree_add_48_2_groupi_n_1016));
 assign csa_tree_add_48_2_groupi_n_1191 = ~((csa_tree_add_48_2_groupi_n_1013 & ~csa_tree_add_48_2_groupi_n_1117)
    | (csa_tree_add_48_2_groupi_n_1014 & csa_tree_add_48_2_groupi_n_1117));
 assign csa_tree_add_48_2_groupi_n_1190 = ~(csa_tree_add_48_2_groupi_n_1150 | csa_tree_add_48_2_groupi_n_41);
 assign csa_tree_add_48_2_groupi_n_1189 = (csa_tree_add_48_2_groupi_n_1113 ^ csa_tree_add_48_2_groupi_n_940);
 assign csa_tree_add_48_2_groupi_n_1185 = ~(csa_tree_add_48_2_groupi_n_1114 ^ csa_tree_add_48_2_groupi_n_942);
 assign csa_tree_add_48_2_groupi_n_1184 = ~csa_tree_add_48_2_groupi_n_1183;
 assign csa_tree_add_48_2_groupi_n_1182 = ~csa_tree_add_48_2_groupi_n_1181;
 assign csa_tree_add_48_2_groupi_n_1179 = ((csa_tree_add_48_2_groupi_n_970 & csa_tree_add_48_2_groupi_n_311)
    | ((csa_tree_add_48_2_groupi_n_311 & csa_tree_add_48_2_groupi_n_998) | (csa_tree_add_48_2_groupi_n_998
    & csa_tree_add_48_2_groupi_n_970)));
 assign csa_tree_add_48_2_groupi_n_1180 = (csa_tree_add_48_2_groupi_n_311 ^ (csa_tree_add_48_2_groupi_n_998
    ^ csa_tree_add_48_2_groupi_n_970));
 assign csa_tree_add_48_2_groupi_n_1177 = ((csa_tree_add_48_2_groupi_n_896 & csa_tree_add_48_2_groupi_n_718)
    | ((csa_tree_add_48_2_groupi_n_718 & csa_tree_add_48_2_groupi_n_965) | (csa_tree_add_48_2_groupi_n_965
    & csa_tree_add_48_2_groupi_n_896)));
 assign csa_tree_add_48_2_groupi_n_1178 = (csa_tree_add_48_2_groupi_n_718 ^ (csa_tree_add_48_2_groupi_n_965
    ^ csa_tree_add_48_2_groupi_n_896));
 assign csa_tree_add_48_2_groupi_n_1175 = ((csa_tree_add_48_2_groupi_n_978 & csa_tree_add_48_2_groupi_n_316)
    | ((csa_tree_add_48_2_groupi_n_316 & csa_tree_add_48_2_groupi_n_720) | (csa_tree_add_48_2_groupi_n_720
    & csa_tree_add_48_2_groupi_n_978)));
 assign csa_tree_add_48_2_groupi_n_1176 = (csa_tree_add_48_2_groupi_n_316 ^ (csa_tree_add_48_2_groupi_n_720
    ^ csa_tree_add_48_2_groupi_n_978));
 assign csa_tree_add_48_2_groupi_n_1181 = ((csa_tree_add_48_2_groupi_n_812 & csa_tree_add_48_2_groupi_n_808)
    | ((csa_tree_add_48_2_groupi_n_808 & csa_tree_add_48_2_groupi_n_807) | (csa_tree_add_48_2_groupi_n_807
    & csa_tree_add_48_2_groupi_n_812)));
 assign csa_tree_add_48_2_groupi_n_1183 = (csa_tree_add_48_2_groupi_n_808 ^ (csa_tree_add_48_2_groupi_n_807
    ^ csa_tree_add_48_2_groupi_n_812));
 assign csa_tree_add_48_2_groupi_n_1173 = ((csa_tree_add_48_2_groupi_n_884 & csa_tree_add_48_2_groupi_n_327)
    | ((csa_tree_add_48_2_groupi_n_327 & csa_tree_add_48_2_groupi_n_919) | (csa_tree_add_48_2_groupi_n_919
    & csa_tree_add_48_2_groupi_n_884)));
 assign csa_tree_add_48_2_groupi_n_1174 = (csa_tree_add_48_2_groupi_n_327 ^ (csa_tree_add_48_2_groupi_n_919
    ^ csa_tree_add_48_2_groupi_n_884));
 assign csa_tree_add_48_2_groupi_n_1171 = ((csa_tree_add_48_2_groupi_n_27 & csa_tree_add_48_2_groupi_n_315)
    | ((csa_tree_add_48_2_groupi_n_315 & csa_tree_add_48_2_groupi_n_322) | (csa_tree_add_48_2_groupi_n_322
    & csa_tree_add_48_2_groupi_n_27)));
 assign csa_tree_add_48_2_groupi_n_1172 = (csa_tree_add_48_2_groupi_n_315 ^ (csa_tree_add_48_2_groupi_n_322
    ^ csa_tree_add_48_2_groupi_n_27));
 assign csa_tree_add_48_2_groupi_n_1169 = ((csa_tree_add_48_2_groupi_n_976 & csa_tree_add_48_2_groupi_n_917)
    | ((csa_tree_add_48_2_groupi_n_917 & csa_tree_add_48_2_groupi_n_25) | (csa_tree_add_48_2_groupi_n_25
    & csa_tree_add_48_2_groupi_n_976)));
 assign csa_tree_add_48_2_groupi_n_1170 = (csa_tree_add_48_2_groupi_n_917 ^ (csa_tree_add_48_2_groupi_n_25
    ^ csa_tree_add_48_2_groupi_n_976));
 assign csa_tree_add_48_2_groupi_n_1167 = ((csa_tree_add_48_2_groupi_n_975 & csa_tree_add_48_2_groupi_n_862)
    | ((csa_tree_add_48_2_groupi_n_862 & csa_tree_add_48_2_groupi_n_717) | (csa_tree_add_48_2_groupi_n_717
    & csa_tree_add_48_2_groupi_n_975)));
 assign csa_tree_add_48_2_groupi_n_1168 = (csa_tree_add_48_2_groupi_n_862 ^ (csa_tree_add_48_2_groupi_n_717
    ^ csa_tree_add_48_2_groupi_n_975));
 assign csa_tree_add_48_2_groupi_n_1165 = ((csa_tree_add_48_2_groupi_n_974 & csa_tree_add_48_2_groupi_n_402)
    | ((csa_tree_add_48_2_groupi_n_402 & csa_tree_add_48_2_groupi_n_715) | (csa_tree_add_48_2_groupi_n_715
    & csa_tree_add_48_2_groupi_n_974)));
 assign csa_tree_add_48_2_groupi_n_1166 = (csa_tree_add_48_2_groupi_n_402 ^ (csa_tree_add_48_2_groupi_n_715
    ^ csa_tree_add_48_2_groupi_n_974));
 assign csa_tree_add_48_2_groupi_n_1163 = ((csa_tree_add_48_2_groupi_n_973 & csa_tree_add_48_2_groupi_n_313)
    | ((csa_tree_add_48_2_groupi_n_313 & csa_tree_add_48_2_groupi_n_719) | (csa_tree_add_48_2_groupi_n_719
    & csa_tree_add_48_2_groupi_n_973)));
 assign csa_tree_add_48_2_groupi_n_1164 = (csa_tree_add_48_2_groupi_n_313 ^ (csa_tree_add_48_2_groupi_n_719
    ^ csa_tree_add_48_2_groupi_n_973));
 assign csa_tree_add_48_2_groupi_n_1161 = ((csa_tree_add_48_2_groupi_n_972 & csa_tree_add_48_2_groupi_n_877)
    | ((csa_tree_add_48_2_groupi_n_877 & csa_tree_add_48_2_groupi_n_716) | (csa_tree_add_48_2_groupi_n_716
    & csa_tree_add_48_2_groupi_n_972)));
 assign csa_tree_add_48_2_groupi_n_1162 = (csa_tree_add_48_2_groupi_n_877 ^ (csa_tree_add_48_2_groupi_n_716
    ^ csa_tree_add_48_2_groupi_n_972));
 assign csa_tree_add_48_2_groupi_n_1160 = ~(csa_tree_add_48_2_groupi_n_1143 & csa_tree_add_48_2_groupi_n_1130);
 assign csa_tree_add_48_2_groupi_n_1159 = ~(csa_tree_add_48_2_groupi_n_1143 | csa_tree_add_48_2_groupi_n_1049);
 assign csa_tree_add_48_2_groupi_n_1158 = ~(csa_tree_add_48_2_groupi_n_1144 | csa_tree_add_48_2_groupi_n_1130);
 assign csa_tree_add_48_2_groupi_n_1157 = ~(csa_tree_add_48_2_groupi_n_1142 | csa_tree_add_48_2_groupi_n_133);
 assign csa_tree_add_48_2_groupi_n_1156 = ~(csa_tree_add_48_2_groupi_n_1142 & csa_tree_add_48_2_groupi_n_133);
 assign csa_tree_add_48_2_groupi_n_1155 = ~(csa_tree_add_48_2_groupi_n_1144 & csa_tree_add_48_2_groupi_n_1049);
 assign csa_tree_add_48_2_groupi_n_1151 = ~(csa_tree_add_48_2_groupi_n_939 & ~(csa_tree_add_48_2_groupi_n_1048
    & csa_tree_add_48_2_groupi_n_406));
 assign csa_tree_add_48_2_groupi_n_1150 = ~(csa_tree_add_48_2_groupi_n_1104 | csa_tree_add_48_2_groupi_n_1014);
 assign csa_tree_add_48_2_groupi_n_1149 = ~(csa_tree_add_48_2_groupi_n_40 | ~csa_tree_add_48_2_groupi_n_1015);
 assign csa_tree_add_48_2_groupi_n_1148 = ~(csa_tree_add_48_2_groupi_n_49 | csa_tree_add_48_2_groupi_n_940);
 assign csa_tree_add_48_2_groupi_n_1147 = ~(csa_tree_add_48_2_groupi_n_1097 | csa_tree_add_48_2_groupi_n_944);
 assign csa_tree_add_48_2_groupi_n_1146 = ~(csa_tree_add_48_2_groupi_n_1096 | csa_tree_add_48_2_groupi_n_942);
 assign csa_tree_add_48_2_groupi_n_1145 = ~(csa_tree_add_48_2_groupi_n_1086 | (csa_tree_add_48_2_groupi_n_1005
    & csa_tree_add_48_2_groupi_n_1073));
 assign csa_tree_add_48_2_groupi_n_1154 = ~(csa_tree_add_48_2_groupi_n_1137 | csa_tree_add_48_2_groupi_n_1139);
 assign csa_tree_add_48_2_groupi_n_1153 = ~(csa_tree_add_48_2_groupi_n_1067 | (csa_tree_add_48_2_groupi_n_1066
    & csa_tree_add_48_2_groupi_n_943));
 assign csa_tree_add_48_2_groupi_n_1152 = ~(csa_tree_add_48_2_groupi_n_1064 & (csa_tree_add_48_2_groupi_n_1062
    | csa_tree_add_48_2_groupi_n_937));
 assign csa_tree_add_48_2_groupi_n_1143 = ~csa_tree_add_48_2_groupi_n_1144;
 assign csa_tree_add_48_2_groupi_n_1142 = ((csa_tree_add_48_2_groupi_n_811 & csa_tree_add_48_2_groupi_n_810)
    | ((csa_tree_add_48_2_groupi_n_810 & csa_tree_add_48_2_groupi_n_809) | (csa_tree_add_48_2_groupi_n_809
    & csa_tree_add_48_2_groupi_n_811)));
 assign csa_tree_add_48_2_groupi_n_1144 = (csa_tree_add_48_2_groupi_n_810 ^ (csa_tree_add_48_2_groupi_n_809
    ^ csa_tree_add_48_2_groupi_n_811));
 assign csa_tree_add_48_2_groupi_n_1140 = (csa_tree_add_48_2_groupi_n_895 & csa_tree_add_48_2_groupi_n_1041);
 assign csa_tree_add_48_2_groupi_n_1141 = (csa_tree_add_48_2_groupi_n_895 ^ csa_tree_add_48_2_groupi_n_1041);
 assign csa_tree_add_48_2_groupi_n_1139 = ~(csa_tree_add_48_2_groupi_n_1126 | csa_tree_add_48_2_groupi_n_1129);
 assign csa_tree_add_48_2_groupi_n_1138 = ~(csa_tree_add_48_2_groupi_n_1126 & csa_tree_add_48_2_groupi_n_1099);
 assign csa_tree_add_48_2_groupi_n_1137 = ~(csa_tree_add_48_2_groupi_n_1125 | csa_tree_add_48_2_groupi_n_1099);
 assign csa_tree_add_48_2_groupi_n_1136 = ~(csa_tree_add_48_2_groupi_n_1125 & csa_tree_add_48_2_groupi_n_1129);
 assign csa_tree_add_48_2_groupi_n_1133 = ~(csa_tree_add_48_2_groupi_n_1091 ^ csa_tree_add_48_2_groupi_n_912);
 assign csa_tree_add_48_2_groupi_n_1135 = ~(csa_tree_add_48_2_groupi_n_988 & (csa_tree_add_48_2_groupi_n_987
    | csa_tree_add_48_2_groupi_n_129));
 assign csa_tree_add_48_2_groupi_n_1132 = ~(csa_tree_add_48_2_groupi_n_1017 ^ (csa_tree_add_48_2_groupi_n_409
    ^ csa_tree_add_48_2_groupi_n_410));
 assign csa_tree_add_48_2_groupi_n_1131 = ~csa_tree_add_48_2_groupi_n_22;
 assign csa_tree_add_48_2_groupi_n_1130 = ~csa_tree_add_48_2_groupi_n_1049;
 assign csa_tree_add_48_2_groupi_n_1129 = ~csa_tree_add_48_2_groupi_n_1099;
 assign csa_tree_add_48_2_groupi_n_1128 = ~n_182;
 assign csa_tree_add_48_2_groupi_n_1127 = ~csa_tree_add_48_2_groupi_n_1046;
 assign csa_tree_add_48_2_groupi_n_1125 = ~csa_tree_add_48_2_groupi_n_1126;
 assign csa_tree_add_48_2_groupi_n_1122 = ((csa_tree_add_48_2_groupi_n_202 & csa_tree_add_48_2_groupi_n_115)
    | ((csa_tree_add_48_2_groupi_n_115 & csa_tree_add_48_2_groupi_n_114) | (csa_tree_add_48_2_groupi_n_114
    & csa_tree_add_48_2_groupi_n_202)));
 assign csa_tree_add_48_2_groupi_n_133 = (csa_tree_add_48_2_groupi_n_115 ^ (csa_tree_add_48_2_groupi_n_114
    ^ csa_tree_add_48_2_groupi_n_202));
 assign csa_tree_add_48_2_groupi_n_1120 = (csa_tree_add_48_2_groupi_n_899 & csa_tree_add_48_2_groupi_n_329);
 assign csa_tree_add_48_2_groupi_n_1121 = (csa_tree_add_48_2_groupi_n_899 ^ csa_tree_add_48_2_groupi_n_329);
 assign csa_tree_add_48_2_groupi_n_1124 = ((csa_tree_add_48_2_groupi_n_684 & csa_tree_add_48_2_groupi_n_683)
    | ((csa_tree_add_48_2_groupi_n_683 & csa_tree_add_48_2_groupi_n_682) | (csa_tree_add_48_2_groupi_n_682
    & csa_tree_add_48_2_groupi_n_684)));
 assign csa_tree_add_48_2_groupi_n_1126 = (csa_tree_add_48_2_groupi_n_683 ^ (csa_tree_add_48_2_groupi_n_682
    ^ csa_tree_add_48_2_groupi_n_684));
 assign csa_tree_add_48_2_groupi_n_1119 = ~((csa_tree_add_48_2_groupi_n_1075 & ~csa_tree_add_48_2_groupi_n_1007)
    | (csa_tree_add_48_2_groupi_n_1074 & csa_tree_add_48_2_groupi_n_1007));
 assign csa_tree_add_48_2_groupi_n_1118 = ~((csa_tree_add_48_2_groupi_n_1081 & ~csa_tree_add_48_2_groupi_n_1002)
    | (csa_tree_add_48_2_groupi_n_1080 & csa_tree_add_48_2_groupi_n_1002));
 assign csa_tree_add_48_2_groupi_n_1117 = ~((csa_tree_add_48_2_groupi_n_1079 & ~csa_tree_add_48_2_groupi_n_1003)
    | (csa_tree_add_48_2_groupi_n_28 & csa_tree_add_48_2_groupi_n_1003));
 assign csa_tree_add_48_2_groupi_n_1114 = ~((csa_tree_add_48_2_groupi_n_1071 & ~csa_tree_add_48_2_groupi_n_1006)
    | (csa_tree_add_48_2_groupi_n_1072 & csa_tree_add_48_2_groupi_n_1006));
 assign csa_tree_add_48_2_groupi_n_1113 = ~((csa_tree_add_48_2_groupi_n_131 & ~csa_tree_add_48_2_groupi_n_130)
    | (csa_tree_add_48_2_groupi_n_1078 & csa_tree_add_48_2_groupi_n_130));
 assign csa_tree_add_48_2_groupi_n_1112 = ~((csa_tree_add_48_2_groupi_n_761 & ~csa_tree_add_48_2_groupi_n_1047)
    | (csa_tree_add_48_2_groupi_n_406 & csa_tree_add_48_2_groupi_n_1047));
 assign csa_tree_add_48_2_groupi_n_1116 = ~(csa_tree_add_48_2_groupi_n_1103 | csa_tree_add_48_2_groupi_n_1101);
 assign csa_tree_add_48_2_groupi_n_1115 = ~(csa_tree_add_48_2_groupi_n_1093 | csa_tree_add_48_2_groupi_n_39);
 assign csa_tree_add_48_2_groupi_n_1111 = ~(csa_tree_add_48_2_groupi_n_1077 & csa_tree_add_48_2_groupi_n_1045);
 assign csa_tree_add_48_2_groupi_n_1110 = ~(csa_tree_add_48_2_groupi_n_1083 | csa_tree_add_48_2_groupi_n_1082);
 assign csa_tree_add_48_2_groupi_n_1109 = ~(csa_tree_add_48_2_groupi_n_1047 & csa_tree_add_48_2_groupi_n_761);
 assign csa_tree_add_48_2_groupi_n_1107 = ~(csa_tree_add_48_2_groupi_n_131 | csa_tree_add_48_2_groupi_n_130);
 assign csa_tree_add_48_2_groupi_n_1106 = ~(csa_tree_add_48_2_groupi_n_1004 & csa_tree_add_48_2_groupi_n_1085);
 assign csa_tree_add_48_2_groupi_n_1105 = ~(csa_tree_add_48_2_groupi_n_1004 | csa_tree_add_48_2_groupi_n_1085);
 assign csa_tree_add_48_2_groupi_n_1104 = ~(csa_tree_add_48_2_groupi_n_1003 | csa_tree_add_48_2_groupi_n_1079);
 assign csa_tree_add_48_2_groupi_n_1103 = ~(csa_tree_add_48_2_groupi_n_1077 | csa_tree_add_48_2_groupi_n_1044);
 assign csa_tree_add_48_2_groupi_n_1102 = ~(csa_tree_add_48_2_groupi_n_1002 | csa_tree_add_48_2_groupi_n_1081);
 assign csa_tree_add_48_2_groupi_n_1101 = ~(csa_tree_add_48_2_groupi_n_1045 | csa_tree_add_48_2_groupi_n_1076);
 assign csa_tree_add_48_2_groupi_n_1100 = ~(csa_tree_add_48_2_groupi_n_1005 | csa_tree_add_48_2_groupi_n_1073);
 assign csa_tree_add_48_2_groupi_n_1097 = ~(csa_tree_add_48_2_groupi_n_1007 | csa_tree_add_48_2_groupi_n_1075);
 assign csa_tree_add_48_2_groupi_n_1096 = ~(csa_tree_add_48_2_groupi_n_1006 | csa_tree_add_48_2_groupi_n_1072);
 assign csa_tree_add_48_2_groupi_n_1095 = ~(csa_tree_add_48_2_groupi_n_1077 | csa_tree_add_48_2_groupi_n_1045);
 assign csa_tree_add_48_2_groupi_n_1094 = ~(csa_tree_add_48_2_groupi_n_1083 & csa_tree_add_48_2_groupi_n_1082);
 assign csa_tree_add_48_2_groupi_n_1093 = ~(csa_tree_add_48_2_groupi_n_1018 | ~(csa_tree_add_48_2_groupi_n_1000
    | csa_tree_add_48_2_groupi_n_750));
 assign csa_tree_add_48_2_groupi_n_1092 = ~((csa_tree_add_48_2_groupi_n_1012 & ~csa_tree_add_48_2_groupi_n_1001)
    | (csa_tree_add_48_2_groupi_n_1011 & csa_tree_add_48_2_groupi_n_1001));
 assign csa_tree_add_48_2_groupi_n_1091 = ~(csa_tree_add_48_2_groupi_n_980 ^ csa_tree_add_48_2_groupi_n_330);
 assign csa_tree_add_48_2_groupi_n_1090 = ~(csa_tree_add_48_2_groupi_n_855 & (csa_tree_add_48_2_groupi_n_1019
    | csa_tree_add_48_2_groupi_n_853));
 assign csa_tree_add_48_2_groupi_n_1099 = ~(csa_tree_add_48_2_groupi_n_713 | (csa_tree_add_48_2_groupi_n_688
    & csa_tree_add_48_2_groupi_n_556));
 assign csa_tree_add_48_2_groupi_n_1089 = (csa_tree_add_48_2_groupi_n_17 ^ csa_tree_add_48_2_groupi_n_556);
 assign csa_tree_add_48_2_groupi_n_1088 = ~(csa_tree_add_48_2_groupi_n_823 & (csa_tree_add_48_2_groupi_n_1017
    | csa_tree_add_48_2_groupi_n_846));
 assign csa_tree_add_48_2_groupi_n_1087 = ~(csa_tree_add_48_2_groupi_n_132 & ~csa_tree_add_48_2_groupi_n_1063);
 assign csa_tree_add_48_2_groupi_n_1085 = ~csa_tree_add_48_2_groupi_n_1084;
 assign csa_tree_add_48_2_groupi_n_1080 = ~csa_tree_add_48_2_groupi_n_1081;
 assign csa_tree_add_48_2_groupi_n_1078 = ~csa_tree_add_48_2_groupi_n_131;
 assign csa_tree_add_48_2_groupi_n_1077 = ~csa_tree_add_48_2_groupi_n_1076;
 assign csa_tree_add_48_2_groupi_n_1074 = ~csa_tree_add_48_2_groupi_n_1075;
 assign csa_tree_add_48_2_groupi_n_1071 = ~csa_tree_add_48_2_groupi_n_1072;
 assign csa_tree_add_48_2_groupi_n_1070 = ~csa_tree_add_48_2_groupi_n_132;
 assign csa_tree_add_48_2_groupi_n_1067 = ~(csa_tree_add_48_2_groupi_n_1012 | csa_tree_add_48_2_groupi_n_1001);
 assign csa_tree_add_48_2_groupi_n_1066 = ~(csa_tree_add_48_2_groupi_n_1012 & csa_tree_add_48_2_groupi_n_1001);
 assign csa_tree_add_48_2_groupi_n_1064 = ~(csa_tree_add_48_2_groupi_n_1009 & csa_tree_add_48_2_groupi_n_1010);
 assign csa_tree_add_48_2_groupi_n_1063 = ~(csa_tree_add_48_2_groupi_n_946 | csa_tree_add_48_2_groupi_n_945);
 assign csa_tree_add_48_2_groupi_n_1062 = ~(csa_tree_add_48_2_groupi_n_1009 | csa_tree_add_48_2_groupi_n_1010);
 assign csa_tree_add_48_2_groupi_n_1061 = ~(csa_tree_add_48_2_groupi_n_758 | (n_185 & {in4[1]}));
 assign csa_tree_add_48_2_groupi_n_1086 = ~(csa_tree_add_48_2_groupi_n_696 | (n_189 & csa_tree_add_48_2_groupi_n_562));
 assign csa_tree_add_48_2_groupi_n_1084 = ~(csa_tree_add_48_2_groupi_n_994 & csa_tree_add_48_2_groupi_n_412);
 assign csa_tree_add_48_2_groupi_n_1060 = ~(csa_tree_add_48_2_groupi_n_412 & (csa_tree_add_48_2_groupi_n_126
    | csa_tree_add_48_2_groupi_n_459));
 assign csa_tree_add_48_2_groupi_n_1059 = ~(csa_tree_add_48_2_groupi_n_304 & (csa_tree_add_48_2_groupi_n_848
    | csa_tree_add_48_2_groupi_n_628));
 assign csa_tree_add_48_2_groupi_n_1058 = ~(csa_tree_add_48_2_groupi_n_754 | (n_189 & {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_1083 = ~(csa_tree_add_48_2_groupi_n_995 | csa_tree_add_48_2_groupi_n_712);
 assign csa_tree_add_48_2_groupi_n_1082 = ~(csa_tree_add_48_2_groupi_n_989 | csa_tree_add_48_2_groupi_n_705);
 assign csa_tree_add_48_2_groupi_n_1081 = ~(csa_tree_add_48_2_groupi_n_6 | csa_tree_add_48_2_groupi_n_693);
 assign csa_tree_add_48_2_groupi_n_1057 = ~(csa_tree_add_48_2_groupi_n_10 & (csa_tree_add_48_2_groupi_n_126
    | csa_tree_add_48_2_groupi_n_460));
 assign csa_tree_add_48_2_groupi_n_1056 = ~(csa_tree_add_48_2_groupi_n_9 & (csa_tree_add_48_2_groupi_n_128
    | csa_tree_add_48_2_groupi_n_480));
 assign csa_tree_add_48_2_groupi_n_1079 = ~(csa_tree_add_48_2_groupi_n_748 & (csa_tree_add_48_2_groupi_n_126
    | csa_tree_add_48_2_groupi_n_487));
 assign csa_tree_add_48_2_groupi_n_1055 = ~(csa_tree_add_48_2_groupi_n_706 & (csa_tree_add_48_2_groupi_n_126
    | csa_tree_add_48_2_groupi_n_457));
 assign csa_tree_add_48_2_groupi_n_131 = ~(csa_tree_add_48_2_groupi_n_992 | csa_tree_add_48_2_groupi_n_710);
 assign csa_tree_add_48_2_groupi_n_1054 = ~(csa_tree_add_48_2_groupi_n_708 & (csa_tree_add_48_2_groupi_n_128
    | csa_tree_add_48_2_groupi_n_476));
 assign csa_tree_add_48_2_groupi_n_1076 = ~(csa_tree_add_48_2_groupi_n_991 | csa_tree_add_48_2_groupi_n_709);
 assign csa_tree_add_48_2_groupi_n_1053 = ~(csa_tree_add_48_2_groupi_n_704 | (n_185 & csa_tree_add_48_2_groupi_n_416));
 assign csa_tree_add_48_2_groupi_n_1075 = ~(csa_tree_add_48_2_groupi_n_711 & (csa_tree_add_48_2_groupi_n_126
    | csa_tree_add_48_2_groupi_n_478));
 assign csa_tree_add_48_2_groupi_n_1073 = ~(csa_tree_add_48_2_groupi_n_990 | csa_tree_add_48_2_groupi_n_707);
 assign csa_tree_add_48_2_groupi_n_1072 = ~(csa_tree_add_48_2_groupi_n_703 & (csa_tree_add_48_2_groupi_n_126
    | csa_tree_add_48_2_groupi_n_490));
 assign csa_tree_add_48_2_groupi_n_1052 = ~(csa_tree_add_48_2_groupi_n_411 & (csa_tree_add_48_2_groupi_n_128
    | csa_tree_add_48_2_groupi_n_489));
 assign csa_tree_add_48_2_groupi_n_132 = ~(csa_tree_add_48_2_groupi_n_946 & csa_tree_add_48_2_groupi_n_945);
 assign csa_tree_add_48_2_groupi_n_1048 = ~csa_tree_add_48_2_groupi_n_1047;
 assign csa_tree_add_48_2_groupi_n_1044 = ~csa_tree_add_48_2_groupi_n_1045;
 assign csa_tree_add_48_2_groupi_n_1043 = ~(csa_tree_add_48_2_groupi_n_985 & csa_tree_add_48_2_groupi_n_691);
 assign csa_tree_add_48_2_groupi_n_1042 = ~(csa_tree_add_48_2_groupi_n_692 | (n_189 & csa_tree_add_48_2_groupi_n_521));
 assign csa_tree_add_48_2_groupi_n_1050 = ~(csa_tree_add_48_2_groupi_n_690 & (csa_tree_add_48_2_groupi_n_848
    | csa_tree_add_48_2_groupi_n_427));
 assign csa_tree_add_48_2_groupi_n_1041 = ~(csa_tree_add_48_2_groupi_n_700 & (csa_tree_add_48_2_groupi_n_848
    | csa_tree_add_48_2_groupi_n_565));
 assign csa_tree_add_48_2_groupi_n_1040 = ~(csa_tree_add_48_2_groupi_n_686 & (csa_tree_add_48_2_groupi_n_848
    | csa_tree_add_48_2_groupi_n_583));
 assign csa_tree_add_48_2_groupi_n_1039 = ~(csa_tree_add_48_2_groupi_n_698 & (csa_tree_add_48_2_groupi_n_848
    | csa_tree_add_48_2_groupi_n_576));
 assign csa_tree_add_48_2_groupi_n_1049 = ~(csa_tree_add_48_2_groupi_n_836 & (csa_tree_add_48_2_groupi_n_837
    | csa_tree_add_48_2_groupi_n_737));
 assign csa_tree_add_48_2_groupi_n_1038 = ~((csa_tree_add_48_2_groupi_n_848 | csa_tree_add_48_2_groupi_n_566)
    & (csa_tree_add_48_2_groupi_n_563 | csa_tree_add_48_2_groupi_n_172));
 assign csa_tree_add_48_2_groupi_n_1037 = ~(csa_tree_add_48_2_groupi_n_986 & csa_tree_add_48_2_groupi_n_685);
 assign csa_tree_add_48_2_groupi_n_1036 = ~(csa_tree_add_48_2_groupi_n_699 & ~(n_189 & csa_tree_add_48_2_groupi_n_572));
 assign csa_tree_add_48_2_groupi_n_130 = ~(csa_tree_add_48_2_groupi_n_697 | (n_189 & csa_tree_add_48_2_groupi_n_569));
 assign csa_tree_add_48_2_groupi_n_1035 = ~(csa_tree_add_48_2_groupi_n_984 & csa_tree_add_48_2_groupi_n_689);
 assign csa_tree_add_48_2_groupi_n_1034 = ~((csa_tree_add_48_2_groupi_n_848 | csa_tree_add_48_2_groupi_n_568)
    & (csa_tree_add_48_2_groupi_n_567 | csa_tree_add_48_2_groupi_n_172));
 assign csa_tree_add_48_2_groupi_n_1033 = ~((csa_tree_add_48_2_groupi_n_848 | csa_tree_add_48_2_groupi_n_557)
    & (csa_tree_add_48_2_groupi_n_566 | csa_tree_add_48_2_groupi_n_172));
 assign csa_tree_add_48_2_groupi_n_1032 = ~((csa_tree_add_48_2_groupi_n_848 | csa_tree_add_48_2_groupi_n_563)
    & (csa_tree_add_48_2_groupi_n_568 | csa_tree_add_48_2_groupi_n_172));
 assign csa_tree_add_48_2_groupi_n_1031 = ~((csa_tree_add_48_2_groupi_n_848 | csa_tree_add_48_2_groupi_n_567)
    & (csa_tree_add_48_2_groupi_n_577 | csa_tree_add_48_2_groupi_n_172));
 assign csa_tree_add_48_2_groupi_n_1047 = ~(csa_tree_add_48_2_groupi_n_694 & (csa_tree_add_48_2_groupi_n_848
    | csa_tree_add_48_2_groupi_n_561));
 assign csa_tree_add_48_2_groupi_n_1030 = ~((csa_tree_add_48_2_groupi_n_848 | csa_tree_add_48_2_groupi_n_611)
    & (csa_tree_add_48_2_groupi_n_612 | csa_tree_add_48_2_groupi_n_172));
 assign csa_tree_add_48_2_groupi_n_1029 = ~(csa_tree_add_48_2_groupi_n_695 & (csa_tree_add_48_2_groupi_n_848
    | csa_tree_add_48_2_groupi_n_575));
 assign csa_tree_add_48_2_groupi_n_1028 = ~((csa_tree_add_48_2_groupi_n_848 | csa_tree_add_48_2_groupi_n_571)
    & (csa_tree_add_48_2_groupi_n_557 | csa_tree_add_48_2_groupi_n_172));
 assign csa_tree_add_48_2_groupi_n_1027 = ~((csa_tree_add_48_2_groupi_n_848 | csa_tree_add_48_2_groupi_n_580)
    & (csa_tree_add_48_2_groupi_n_559 | csa_tree_add_48_2_groupi_n_172));
 assign csa_tree_add_48_2_groupi_n_1026 = ~((csa_tree_add_48_2_groupi_n_848 | csa_tree_add_48_2_groupi_n_578)
    & (csa_tree_add_48_2_groupi_n_611 | csa_tree_add_48_2_groupi_n_172));
 assign csa_tree_add_48_2_groupi_n_1025 = ~((csa_tree_add_48_2_groupi_n_848 | csa_tree_add_48_2_groupi_n_559)
    & (csa_tree_add_48_2_groupi_n_571 | csa_tree_add_48_2_groupi_n_172));
 assign csa_tree_add_48_2_groupi_n_1024 = ~((csa_tree_add_48_2_groupi_n_848 | csa_tree_add_48_2_groupi_n_612)
    & (csa_tree_add_48_2_groupi_n_629 | csa_tree_add_48_2_groupi_n_172));
 assign csa_tree_add_48_2_groupi_n_1023 = ~((csa_tree_add_48_2_groupi_n_848 | csa_tree_add_48_2_groupi_n_629)
    & (csa_tree_add_48_2_groupi_n_627 | csa_tree_add_48_2_groupi_n_172));
 assign csa_tree_add_48_2_groupi_n_1022 = ~((csa_tree_add_48_2_groupi_n_848 | csa_tree_add_48_2_groupi_n_627)
    & (csa_tree_add_48_2_groupi_n_628 | csa_tree_add_48_2_groupi_n_172));
 assign csa_tree_add_48_2_groupi_n_1021 = ~((csa_tree_add_48_2_groupi_n_848 | csa_tree_add_48_2_groupi_n_577)
    & (csa_tree_add_48_2_groupi_n_578 | csa_tree_add_48_2_groupi_n_172));
 assign csa_tree_add_48_2_groupi_n_1046 = ~(csa_tree_add_48_2_groupi_n_983 | csa_tree_add_48_2_groupi_n_838);
 assign csa_tree_add_48_2_groupi_n_1045 = ~(csa_tree_add_48_2_groupi_n_18 & csa_tree_add_48_2_groupi_n_687);
 assign csa_tree_add_48_2_groupi_n_1014 = ~csa_tree_add_48_2_groupi_n_1013;
 assign csa_tree_add_48_2_groupi_n_1012 = ~csa_tree_add_48_2_groupi_n_1011;
 assign csa_tree_add_48_2_groupi_n_1009 = ~csa_tree_add_48_2_groupi_n_1008;
 assign csa_tree_add_48_2_groupi_n_999 = ~csa_tree_add_48_2_groupi_n_998;
 assign csa_tree_add_48_2_groupi_n_997 = ~csa_tree_add_48_2_groupi_n_996;
 assign csa_tree_add_48_2_groupi_n_995 = ~(csa_tree_add_48_2_groupi_n_128 | csa_tree_add_48_2_groupi_n_430);
 assign csa_tree_add_48_2_groupi_n_994 = ~(n_187 & {in6[1]});
 assign csa_tree_add_48_2_groupi_n_993 = ~(csa_tree_add_48_2_groupi_n_126 | csa_tree_add_48_2_groupi_n_487);
 assign csa_tree_add_48_2_groupi_n_992 = ~(csa_tree_add_48_2_groupi_n_128 | csa_tree_add_48_2_groupi_n_472);
 assign csa_tree_add_48_2_groupi_n_991 = ~(csa_tree_add_48_2_groupi_n_128 | csa_tree_add_48_2_groupi_n_451);
 assign csa_tree_add_48_2_groupi_n_990 = (n_185 & csa_tree_add_48_2_groupi_n_471);
 assign csa_tree_add_48_2_groupi_n_989 = ~(csa_tree_add_48_2_groupi_n_126 | csa_tree_add_48_2_groupi_n_422);
 assign csa_tree_add_48_2_groupi_n_988 = ~(csa_tree_add_48_2_groupi_n_850 & csa_tree_add_48_2_groupi_n_851);
 assign csa_tree_add_48_2_groupi_n_987 = ~(csa_tree_add_48_2_groupi_n_850 | csa_tree_add_48_2_groupi_n_851);
 assign csa_tree_add_48_2_groupi_n_986 = ~(n_189 & csa_tree_add_48_2_groupi_n_581);
 assign csa_tree_add_48_2_groupi_n_985 = ~(n_189 & csa_tree_add_48_2_groupi_n_573);
 assign csa_tree_add_48_2_groupi_n_984 = ~(n_189 & csa_tree_add_48_2_groupi_n_570);
 assign csa_tree_add_48_2_groupi_n_983 = ~(csa_tree_add_48_2_groupi_n_739 | (csa_tree_add_48_2_groupi_n_733
    & csa_tree_add_48_2_groupi_n_734));
 assign csa_tree_add_48_2_groupi_n_982 = ~((csa_tree_add_48_2_groupi_n_739 & ~csa_tree_add_48_2_groupi_n_732)
    | (csa_tree_add_48_2_groupi_n_738 & csa_tree_add_48_2_groupi_n_732));
 assign csa_tree_add_48_2_groupi_n_981 = ~((csa_tree_add_48_2_groupi_n_737 & ~csa_tree_add_48_2_groupi_n_735)
    | (csa_tree_add_48_2_groupi_n_736 & csa_tree_add_48_2_groupi_n_735));
 assign csa_tree_add_48_2_groupi_n_980 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_622)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_171));
 assign csa_tree_add_48_2_groupi_n_979 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_632)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_530));
 assign csa_tree_add_48_2_groupi_n_1020 = ~(csa_tree_add_48_2_groupi_n_852 & ~csa_tree_add_48_2_groupi_n_854);
 assign csa_tree_add_48_2_groupi_n_978 = ~(csa_tree_add_48_2_groupi_n_788 & csa_tree_add_48_2_groupi_n_825);
 assign csa_tree_add_48_2_groupi_n_977 = ~(csa_tree_add_48_2_groupi_n_786 & csa_tree_add_48_2_groupi_n_820);
 assign csa_tree_add_48_2_groupi_n_976 = ~(csa_tree_add_48_2_groupi_n_795 & csa_tree_add_48_2_groupi_n_816);
 assign csa_tree_add_48_2_groupi_n_1019 = ~(csa_tree_add_48_2_groupi_n_29 | csa_tree_add_48_2_groupi_n_818);
 assign csa_tree_add_48_2_groupi_n_975 = ~(csa_tree_add_48_2_groupi_n_743 | (csa_tree_add_48_2_groupi_n_724
    & {in4[7]}));
 assign csa_tree_add_48_2_groupi_n_974 = ~(csa_tree_add_48_2_groupi_n_741 | (csa_tree_add_48_2_groupi_n_125
    & {in6[7]}));
 assign csa_tree_add_48_2_groupi_n_973 = ~(csa_tree_add_48_2_groupi_n_790 & csa_tree_add_48_2_groupi_n_742);
 assign csa_tree_add_48_2_groupi_n_972 = ~(csa_tree_add_48_2_groupi_n_793 & csa_tree_add_48_2_groupi_n_740);
 assign csa_tree_add_48_2_groupi_n_1018 = ~(csa_tree_add_48_2_groupi_n_785 | csa_tree_add_48_2_groupi_n_30);
 assign csa_tree_add_48_2_groupi_n_1017 = ~(csa_tree_add_48_2_groupi_n_789 | csa_tree_add_48_2_groupi_n_819);
 assign csa_tree_add_48_2_groupi_n_971 = ~(csa_tree_add_48_2_groupi_n_798 & csa_tree_add_48_2_groupi_n_656);
 assign csa_tree_add_48_2_groupi_n_1016 = ~(csa_tree_add_48_2_groupi_n_8 | csa_tree_add_48_2_groupi_n_5);
 assign csa_tree_add_48_2_groupi_n_970 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_607)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_632));
 assign csa_tree_add_48_2_groupi_n_969 = ~(csa_tree_add_48_2_groupi_n_839 & csa_tree_add_48_2_groupi_n_676);
 assign csa_tree_add_48_2_groupi_n_968 = ~(csa_tree_add_48_2_groupi_n_800 & csa_tree_add_48_2_groupi_n_671);
 assign csa_tree_add_48_2_groupi_n_967 = ~(csa_tree_add_48_2_groupi_n_814 & csa_tree_add_48_2_groupi_n_665);
 assign csa_tree_add_48_2_groupi_n_966 = ~(csa_tree_add_48_2_groupi_n_842 & csa_tree_add_48_2_groupi_n_666);
 assign csa_tree_add_48_2_groupi_n_1015 = ~(csa_tree_add_48_2_groupi_n_804 & csa_tree_add_48_2_groupi_n_677);
 assign csa_tree_add_48_2_groupi_n_1013 = ~(csa_tree_add_48_2_groupi_n_834 & csa_tree_add_48_2_groupi_n_669);
 assign csa_tree_add_48_2_groupi_n_965 = ~(csa_tree_add_48_2_groupi_n_831 | csa_tree_add_48_2_groupi_n_747);
 assign csa_tree_add_48_2_groupi_n_964 = ~(csa_tree_add_48_2_groupi_n_3 | csa_tree_add_48_2_groupi_n_670);
 assign csa_tree_add_48_2_groupi_n_963 = ~(csa_tree_add_48_2_groupi_n_845 | csa_tree_add_48_2_groupi_n_673);
 assign csa_tree_add_48_2_groupi_n_962 = ~(csa_tree_add_48_2_groupi_n_833 & csa_tree_add_48_2_groupi_n_658);
 assign csa_tree_add_48_2_groupi_n_961 = ~(csa_tree_add_48_2_groupi_n_841 & csa_tree_add_48_2_groupi_n_654);
 assign csa_tree_add_48_2_groupi_n_960 = ~(csa_tree_add_48_2_groupi_n_7 & csa_tree_add_48_2_groupi_n_664);
 assign csa_tree_add_48_2_groupi_n_959 = ~(csa_tree_add_48_2_groupi_n_702 & ~(csa_tree_add_48_2_groupi_n_721
    & csa_tree_add_48_2_groupi_n_449));
 assign csa_tree_add_48_2_groupi_n_1011 = ~(csa_tree_add_48_2_groupi_n_829 & csa_tree_add_48_2_groupi_n_668);
 assign csa_tree_add_48_2_groupi_n_1010 = ~(csa_tree_add_48_2_groupi_n_803 & csa_tree_add_48_2_groupi_n_659);
 assign csa_tree_add_48_2_groupi_n_1008 = ~(csa_tree_add_48_2_groupi_n_675 | ~(csa_tree_add_48_2_groupi_n_722
    | csa_tree_add_48_2_groupi_n_461));
 assign csa_tree_add_48_2_groupi_n_958 = ~(csa_tree_add_48_2_groupi_n_840 & csa_tree_add_48_2_groupi_n_662);
 assign csa_tree_add_48_2_groupi_n_1007 = ~(csa_tree_add_48_2_groupi_n_843 & csa_tree_add_48_2_groupi_n_4);
 assign csa_tree_add_48_2_groupi_n_1006 = ~(csa_tree_add_48_2_groupi_n_781 & csa_tree_add_48_2_groupi_n_672);
 assign csa_tree_add_48_2_groupi_n_1005 = ~(csa_tree_add_48_2_groupi_n_805 | csa_tree_add_48_2_groupi_n_660);
 assign csa_tree_add_48_2_groupi_n_1004 = ~(csa_tree_add_48_2_groupi_n_828 & csa_tree_add_48_2_groupi_n_674);
 assign csa_tree_add_48_2_groupi_n_957 = ~(csa_tree_add_48_2_groupi_n_801 & csa_tree_add_48_2_groupi_n_661);
 assign csa_tree_add_48_2_groupi_n_956 = ~(csa_tree_add_48_2_groupi_n_815 & csa_tree_add_48_2_groupi_n_701);
 assign csa_tree_add_48_2_groupi_n_1003 = ~(csa_tree_add_48_2_groupi_n_832 & csa_tree_add_48_2_groupi_n_667);
 assign csa_tree_add_48_2_groupi_n_1002 = ~(csa_tree_add_48_2_groupi_n_16 | ~(csa_tree_add_48_2_groupi_n_726
    | csa_tree_add_48_2_groupi_n_466));
 assign csa_tree_add_48_2_groupi_n_955 = ~(csa_tree_add_48_2_groupi_n_813 & csa_tree_add_48_2_groupi_n_657);
 assign csa_tree_add_48_2_groupi_n_954 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_618)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_622));
 assign csa_tree_add_48_2_groupi_n_953 = ~(csa_tree_add_48_2_groupi_n_663 & ~(csa_tree_add_48_2_groupi_n_721
    & csa_tree_add_48_2_groupi_n_447));
 assign csa_tree_add_48_2_groupi_n_952 = ~(csa_tree_add_48_2_groupi_n_21 | csa_tree_add_48_2_groupi_n_745);
 assign csa_tree_add_48_2_groupi_n_1001 = ~(csa_tree_add_48_2_groupi_n_794 | csa_tree_add_48_2_groupi_n_822);
 assign csa_tree_add_48_2_groupi_n_1000 = ~(csa_tree_add_48_2_groupi_n_799 & csa_tree_add_48_2_groupi_n_746);
 assign csa_tree_add_48_2_groupi_n_951 = ~(csa_tree_add_48_2_groupi_n_835 & csa_tree_add_48_2_groupi_n_744);
 assign csa_tree_add_48_2_groupi_n_950 = ~(csa_tree_add_48_2_groupi_n_784 & csa_tree_add_48_2_groupi_n_821);
 assign csa_tree_add_48_2_groupi_n_949 = ~(csa_tree_add_48_2_groupi_n_787 & csa_tree_add_48_2_groupi_n_824);
 assign csa_tree_add_48_2_groupi_n_948 = ~(csa_tree_add_48_2_groupi_n_792 | csa_tree_add_48_2_groupi_n_847);
 assign csa_tree_add_48_2_groupi_n_947 = ~(csa_tree_add_48_2_groupi_n_791 & ~(csa_tree_add_48_2_groupi_n_550
    & csa_tree_add_48_2_groupi_n_752));
 assign csa_tree_add_48_2_groupi_n_998 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_613)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_618));
 assign csa_tree_add_48_2_groupi_n_996 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_609)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_613));
 assign csa_tree_add_48_2_groupi_n_939 = ~csa_tree_add_48_2_groupi_n_938;
 assign csa_tree_add_48_2_groupi_n_936 = ~csa_tree_add_48_2_groupi_n_935;
 assign csa_tree_add_48_2_groupi_n_934 = ~csa_tree_add_48_2_groupi_n_933;
 assign csa_tree_add_48_2_groupi_n_932 = ~csa_tree_add_48_2_groupi_n_931;
 assign csa_tree_add_48_2_groupi_n_930 = ~csa_tree_add_48_2_groupi_n_929;
 assign csa_tree_add_48_2_groupi_n_928 = ~csa_tree_add_48_2_groupi_n_927;
 assign csa_tree_add_48_2_groupi_n_926 = ~csa_tree_add_48_2_groupi_n_925;
 assign csa_tree_add_48_2_groupi_n_924 = ~csa_tree_add_48_2_groupi_n_923;
 assign csa_tree_add_48_2_groupi_n_922 = ~csa_tree_add_48_2_groupi_n_921;
 assign csa_tree_add_48_2_groupi_n_920 = ~csa_tree_add_48_2_groupi_n_919;
 assign csa_tree_add_48_2_groupi_n_918 = ~csa_tree_add_48_2_groupi_n_917;
 assign csa_tree_add_48_2_groupi_n_916 = ~csa_tree_add_48_2_groupi_n_915;
 assign csa_tree_add_48_2_groupi_n_914 = ~csa_tree_add_48_2_groupi_n_913;
 assign csa_tree_add_48_2_groupi_n_946 = ~(csa_tree_add_48_2_groupi_n_645 | ~(csa_tree_add_48_2_groupi_n_122
    | csa_tree_add_48_2_groupi_n_616));
 assign csa_tree_add_48_2_groupi_n_912 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_614)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_523));
 assign csa_tree_add_48_2_groupi_n_945 = ~(csa_tree_add_48_2_groupi_n_777 | ~(csa_tree_add_48_2_groupi_n_680
    | csa_tree_add_48_2_groupi_n_762));
 assign csa_tree_add_48_2_groupi_n_911 = ~(csa_tree_add_48_2_groupi_n_765 & csa_tree_add_48_2_groupi_n_778);
 assign csa_tree_add_48_2_groupi_n_910 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_499)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_519));
 assign csa_tree_add_48_2_groupi_n_944 = ~(csa_tree_add_48_2_groupi_n_1 | csa_tree_add_48_2_groupi_n_2);
 assign csa_tree_add_48_2_groupi_n_943 = ~(csa_tree_add_48_2_groupi_n_764 & csa_tree_add_48_2_groupi_n_780);
 assign csa_tree_add_48_2_groupi_n_942 = ~(csa_tree_add_48_2_groupi_n_766 | csa_tree_add_48_2_groupi_n_635);
 assign csa_tree_add_48_2_groupi_n_909 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_601)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_614));
 assign csa_tree_add_48_2_groupi_n_908 = ~(csa_tree_add_48_2_groupi_n_771 & csa_tree_add_48_2_groupi_n_639);
 assign csa_tree_add_48_2_groupi_n_907 = ~(csa_tree_add_48_2_groupi_n_19 & csa_tree_add_48_2_groupi_n_643);
 assign csa_tree_add_48_2_groupi_n_941 = ~(csa_tree_add_48_2_groupi_n_770 | csa_tree_add_48_2_groupi_n_641);
 assign csa_tree_add_48_2_groupi_n_940 = ~(csa_tree_add_48_2_groupi_n_20 | csa_tree_add_48_2_groupi_n_642);
 assign csa_tree_add_48_2_groupi_n_906 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_626)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_431));
 assign csa_tree_add_48_2_groupi_n_905 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_431)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_440));
 assign csa_tree_add_48_2_groupi_n_904 = ~(csa_tree_add_48_2_groupi_n_15 & csa_tree_add_48_2_groupi_n_648);
 assign csa_tree_add_48_2_groupi_n_903 = ~(csa_tree_add_48_2_groupi_n_779 & ~(csa_tree_add_48_2_groupi_n_681
    & csa_tree_add_48_2_groupi_n_596));
 assign csa_tree_add_48_2_groupi_n_902 = ~(csa_tree_add_48_2_groupi_n_31 & csa_tree_add_48_2_groupi_n_806);
 assign csa_tree_add_48_2_groupi_n_901 = ~(csa_tree_add_48_2_groupi_n_782 & ~(csa_tree_add_48_2_groupi_n_681
    & csa_tree_add_48_2_groupi_n_603));
 assign csa_tree_add_48_2_groupi_n_900 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_589)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_587));
 assign csa_tree_add_48_2_groupi_n_899 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_516)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_500));
 assign csa_tree_add_48_2_groupi_n_898 = ~(csa_tree_add_48_2_groupi_n_767 & csa_tree_add_48_2_groupi_n_636);
 assign csa_tree_add_48_2_groupi_n_897 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_507)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_520));
 assign csa_tree_add_48_2_groupi_n_896 = ~(csa_tree_add_48_2_groupi_n_776 & ~(csa_tree_add_48_2_groupi_n_681
    & csa_tree_add_48_2_groupi_n_591));
 assign csa_tree_add_48_2_groupi_n_895 = ~(csa_tree_add_48_2_groupi_n_650 & ~(csa_tree_add_48_2_groupi_n_123
    & csa_tree_add_48_2_groupi_n_510));
 assign csa_tree_add_48_2_groupi_n_894 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_504)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_502));
 assign csa_tree_add_48_2_groupi_n_893 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_503)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_499));
 assign csa_tree_add_48_2_groupi_n_892 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_513)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_509));
 assign csa_tree_add_48_2_groupi_n_891 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_520)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_506));
 assign csa_tree_add_48_2_groupi_n_890 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_502)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_507));
 assign csa_tree_add_48_2_groupi_n_889 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_509)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_504));
 assign csa_tree_add_48_2_groupi_n_938 = ~(csa_tree_add_48_2_groupi_n_13 | csa_tree_add_48_2_groupi_n_14);
 assign csa_tree_add_48_2_groupi_n_888 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_498)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_516));
 assign csa_tree_add_48_2_groupi_n_887 = ~(csa_tree_add_48_2_groupi_n_647 | ~(csa_tree_add_48_2_groupi_n_679
    | csa_tree_add_48_2_groupi_n_508));
 assign csa_tree_add_48_2_groupi_n_886 = ~(csa_tree_add_48_2_groupi_n_774 & csa_tree_add_48_2_groupi_n_652);
 assign csa_tree_add_48_2_groupi_n_885 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_608)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_607));
 assign csa_tree_add_48_2_groupi_n_884 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_501)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_503));
 assign csa_tree_add_48_2_groupi_n_883 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_506)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_608));
 assign csa_tree_add_48_2_groupi_n_882 = ~(csa_tree_add_48_2_groupi_n_646 & ~(csa_tree_add_48_2_groupi_n_123
    & csa_tree_add_48_2_groupi_n_512));
 assign csa_tree_add_48_2_groupi_n_881 = ~(csa_tree_add_48_2_groupi_n_773 & csa_tree_add_48_2_groupi_n_11);
 assign csa_tree_add_48_2_groupi_n_880 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_519)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_513));
 assign csa_tree_add_48_2_groupi_n_937 = ~(csa_tree_add_48_2_groupi_n_772 | csa_tree_add_48_2_groupi_n_12);
 assign csa_tree_add_48_2_groupi_n_879 = ~(csa_tree_add_48_2_groupi_n_651 & ~(csa_tree_add_48_2_groupi_n_123
    & csa_tree_add_48_2_groupi_n_517));
 assign csa_tree_add_48_2_groupi_n_878 = ~(csa_tree_add_48_2_groupi_n_797 & csa_tree_add_48_2_groupi_n_827);
 assign csa_tree_add_48_2_groupi_n_877 = ~(csa_tree_add_48_2_groupi_n_649 & ~(csa_tree_add_48_2_groupi_n_123
    & csa_tree_add_48_2_groupi_n_505));
 assign csa_tree_add_48_2_groupi_n_876 = ~((csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_500)
    & (csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_501));
 assign csa_tree_add_48_2_groupi_n_875 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_590)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_602));
 assign csa_tree_add_48_2_groupi_n_874 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_586)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_599));
 assign csa_tree_add_48_2_groupi_n_873 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_599)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_606));
 assign csa_tree_add_48_2_groupi_n_872 = ~(csa_tree_add_48_2_groupi_n_763 & csa_tree_add_48_2_groupi_n_775);
 assign csa_tree_add_48_2_groupi_n_871 = ~(csa_tree_add_48_2_groupi_n_796 & csa_tree_add_48_2_groupi_n_826);
 assign csa_tree_add_48_2_groupi_n_870 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_587)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_595));
 assign csa_tree_add_48_2_groupi_n_869 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_631)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_626));
 assign csa_tree_add_48_2_groupi_n_868 = ~(csa_tree_add_48_2_groupi_n_768 & csa_tree_add_48_2_groupi_n_638);
 assign csa_tree_add_48_2_groupi_n_867 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_606)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_601));
 assign csa_tree_add_48_2_groupi_n_866 = ~(csa_tree_add_48_2_groupi_n_769 & csa_tree_add_48_2_groupi_n_644);
 assign csa_tree_add_48_2_groupi_n_865 = ~(csa_tree_add_48_2_groupi_n_783 & csa_tree_add_48_2_groupi_n_817);
 assign csa_tree_add_48_2_groupi_n_864 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_440)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_435));
 assign csa_tree_add_48_2_groupi_n_863 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_592)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_593));
 assign csa_tree_add_48_2_groupi_n_862 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_760)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_590));
 assign csa_tree_add_48_2_groupi_n_861 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_595)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_585));
 assign csa_tree_add_48_2_groupi_n_860 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_594)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_588));
 assign csa_tree_add_48_2_groupi_n_859 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_593)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_586));
 assign csa_tree_add_48_2_groupi_n_858 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_597)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_594));
 assign csa_tree_add_48_2_groupi_n_857 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_588)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_592));
 assign csa_tree_add_48_2_groupi_n_856 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_585)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_597));
 assign csa_tree_add_48_2_groupi_n_935 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_619)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_436));
 assign csa_tree_add_48_2_groupi_n_933 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_621)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_610));
 assign csa_tree_add_48_2_groupi_n_931 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_436)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_433));
 assign csa_tree_add_48_2_groupi_n_929 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_439)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_619));
 assign csa_tree_add_48_2_groupi_n_927 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_438)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_439));
 assign csa_tree_add_48_2_groupi_n_925 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_432)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_438));
 assign csa_tree_add_48_2_groupi_n_923 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_433)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_621));
 assign csa_tree_add_48_2_groupi_n_921 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_610)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_609));
 assign csa_tree_add_48_2_groupi_n_919 = ~((csa_tree_add_48_2_groupi_n_680 | csa_tree_add_48_2_groupi_n_602)
    & (csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_589));
 assign csa_tree_add_48_2_groupi_n_917 = ~(csa_tree_add_48_2_groupi_n_640 & ~(csa_tree_add_48_2_groupi_n_121
    & csa_tree_add_48_2_groupi_n_625));
 assign csa_tree_add_48_2_groupi_n_915 = ~(csa_tree_add_48_2_groupi_n_0 | csa_tree_add_48_2_groupi_n_637);
 assign csa_tree_add_48_2_groupi_n_913 = ~((csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_435)
    & (csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_432));
 assign csa_tree_add_48_2_groupi_n_855 = ~csa_tree_add_48_2_groupi_n_854;
 assign csa_tree_add_48_2_groupi_n_853 = ~csa_tree_add_48_2_groupi_n_852;
 assign csa_tree_add_48_2_groupi_n_128 = ~n_185;
 assign csa_tree_add_48_2_groupi_n_126 = ~n_187;
 assign csa_tree_add_48_2_groupi_n_848 = ~n_189;
 assign csa_tree_add_48_2_groupi_n_847 = ~(csa_tree_add_48_2_groupi_n_553 | csa_tree_add_48_2_groupi_n_491);
 assign csa_tree_add_48_2_groupi_n_846 = (csa_tree_add_48_2_groupi_n_409 & csa_tree_add_48_2_groupi_n_410);
 assign csa_tree_add_48_2_groupi_n_845 = ~(csa_tree_add_48_2_groupi_n_722 | csa_tree_add_48_2_groupi_n_455);
 assign csa_tree_add_48_2_groupi_n_844 = ~(csa_tree_add_48_2_groupi_n_730 & csa_tree_add_48_2_groupi_n_456);
 assign csa_tree_add_48_2_groupi_n_843 = ~(csa_tree_add_48_2_groupi_n_727 & csa_tree_add_48_2_groupi_n_463);
 assign csa_tree_add_48_2_groupi_n_842 = ~(csa_tree_add_48_2_groupi_n_730 & csa_tree_add_48_2_groupi_n_473);
 assign csa_tree_add_48_2_groupi_n_841 = ~(csa_tree_add_48_2_groupi_n_721 & ~csa_tree_add_48_2_groupi_n_464);
 assign csa_tree_add_48_2_groupi_n_840 = ~(csa_tree_add_48_2_groupi_n_728 & csa_tree_add_48_2_groupi_n_454);
 assign csa_tree_add_48_2_groupi_n_839 = ~(csa_tree_add_48_2_groupi_n_728 & csa_tree_add_48_2_groupi_n_453);
 assign csa_tree_add_48_2_groupi_n_838 = ~(csa_tree_add_48_2_groupi_n_733 | csa_tree_add_48_2_groupi_n_734);
 assign csa_tree_add_48_2_groupi_n_837 = ~(csa_tree_add_48_2_groupi_n_735 | csa_tree_add_48_2_groupi_n_731);
 assign csa_tree_add_48_2_groupi_n_836 = ~(csa_tree_add_48_2_groupi_n_735 & csa_tree_add_48_2_groupi_n_731);
 assign csa_tree_add_48_2_groupi_n_835 = ~(csa_tree_add_48_2_groupi_n_727 & csa_tree_add_48_2_groupi_n_450);
 assign csa_tree_add_48_2_groupi_n_834 = ~(csa_tree_add_48_2_groupi_n_730 & csa_tree_add_48_2_groupi_n_479);
 assign csa_tree_add_48_2_groupi_n_833 = ~(csa_tree_add_48_2_groupi_n_728 & csa_tree_add_48_2_groupi_n_488);
 assign csa_tree_add_48_2_groupi_n_832 = ~(csa_tree_add_48_2_groupi_n_727 & csa_tree_add_48_2_groupi_n_485);
 assign csa_tree_add_48_2_groupi_n_831 = ~(csa_tree_add_48_2_groupi_n_729 | csa_tree_add_48_2_groupi_n_174);
 assign csa_tree_add_48_2_groupi_n_830 = ~(csa_tree_add_48_2_groupi_n_722 | csa_tree_add_48_2_groupi_n_175);
 assign csa_tree_add_48_2_groupi_n_829 = ~(csa_tree_add_48_2_groupi_n_728 & csa_tree_add_48_2_groupi_n_469);
 assign csa_tree_add_48_2_groupi_n_828 = ~(csa_tree_add_48_2_groupi_n_727 & csa_tree_add_48_2_groupi_n_484);
 assign csa_tree_add_48_2_groupi_n_827 = ~(csa_tree_add_48_2_groupi_n_552 & csa_tree_add_48_2_groupi_n_493);
 assign csa_tree_add_48_2_groupi_n_826 = ~(csa_tree_add_48_2_groupi_n_550 & csa_tree_add_48_2_groupi_n_494);
 assign csa_tree_add_48_2_groupi_n_825 = ~(csa_tree_add_48_2_groupi_n_552 & csa_tree_add_48_2_groupi_n_755);
 assign csa_tree_add_48_2_groupi_n_824 = ~(csa_tree_add_48_2_groupi_n_550 & csa_tree_add_48_2_groupi_n_756);
 assign csa_tree_add_48_2_groupi_n_823 = (csa_tree_add_48_2_groupi_n_409 | csa_tree_add_48_2_groupi_n_410);
 assign csa_tree_add_48_2_groupi_n_822 = ~(csa_tree_add_48_2_groupi_n_549 | csa_tree_add_48_2_groupi_n_497);
 assign csa_tree_add_48_2_groupi_n_821 = ~(csa_tree_add_48_2_groupi_n_552 & csa_tree_add_48_2_groupi_n_757);
 assign csa_tree_add_48_2_groupi_n_820 = ~(csa_tree_add_48_2_groupi_n_552 & csa_tree_add_48_2_groupi_n_759);
 assign csa_tree_add_48_2_groupi_n_819 = ~(csa_tree_add_48_2_groupi_n_549 | csa_tree_add_48_2_groupi_n_496);
 assign csa_tree_add_48_2_groupi_n_818 = ~(csa_tree_add_48_2_groupi_n_549 | csa_tree_add_48_2_groupi_n_495);
 assign csa_tree_add_48_2_groupi_n_817 = ~(csa_tree_add_48_2_groupi_n_552 & csa_tree_add_48_2_groupi_n_492);
 assign csa_tree_add_48_2_groupi_n_816 = ~(csa_tree_add_48_2_groupi_n_550 & csa_tree_add_48_2_groupi_n_753);
 assign csa_tree_add_48_2_groupi_n_815 = ~(csa_tree_add_48_2_groupi_n_727 & csa_tree_add_48_2_groupi_n_462);
 assign csa_tree_add_48_2_groupi_n_814 = ~(csa_tree_add_48_2_groupi_n_730 & csa_tree_add_48_2_groupi_n_475);
 assign csa_tree_add_48_2_groupi_n_813 = ~(csa_tree_add_48_2_groupi_n_728 & csa_tree_add_48_2_groupi_n_483);
 assign csa_tree_add_48_2_groupi_n_854 = ~(csa_tree_add_48_2_groupi_n_414 | csa_tree_add_48_2_groupi_n_413);
 assign csa_tree_add_48_2_groupi_n_852 = ~(csa_tree_add_48_2_groupi_n_414 & csa_tree_add_48_2_groupi_n_413);
 assign csa_tree_add_48_2_groupi_n_812 = ~(csa_tree_add_48_2_groupi_n_655 & {in2[5]});
 assign csa_tree_add_48_2_groupi_n_811 = ~(csa_tree_add_48_2_groupi_n_173 | (csa_tree_add_48_2_groupi_n_540
    & csa_tree_add_48_2_groupi_n_110));
 assign csa_tree_add_48_2_groupi_n_129 = ~({in2[3]} & (csa_tree_add_48_2_groupi_n_533 | csa_tree_add_48_2_groupi_n_395));
 assign csa_tree_add_48_2_groupi_n_810 = ~(csa_tree_add_48_2_groupi_n_136 | (csa_tree_add_48_2_groupi_n_535
    & csa_tree_add_48_2_groupi_n_112));
 assign csa_tree_add_48_2_groupi_n_851 = ~(csa_tree_add_48_2_groupi_n_653 | csa_tree_add_48_2_groupi_n_175);
 assign csa_tree_add_48_2_groupi_n_809 = ~(csa_tree_add_48_2_groupi_n_139 | (csa_tree_add_48_2_groupi_n_539
    & csa_tree_add_48_2_groupi_n_113));
 assign csa_tree_add_48_2_groupi_n_850 = ~(csa_tree_add_48_2_groupi_n_634 | csa_tree_add_48_2_groupi_n_140);
 assign csa_tree_add_48_2_groupi_n_808 = ~({in6[5]} & (csa_tree_add_48_2_groupi_n_522 | csa_tree_add_48_2_groupi_n_399));
 assign csa_tree_add_48_2_groupi_n_807 = ~({in4[5]} & (csa_tree_add_48_2_groupi_n_538 | csa_tree_add_48_2_groupi_n_400));
 assign csa_tree_add_48_2_groupi_n_806 = ~(csa_tree_add_48_2_groupi_n_546 & csa_tree_add_48_2_groupi_n_603);
 assign csa_tree_add_48_2_groupi_n_805 = (csa_tree_add_48_2_groupi_n_721 & csa_tree_add_48_2_groupi_n_421);
 assign csa_tree_add_48_2_groupi_n_804 = ~(csa_tree_add_48_2_groupi_n_730 & csa_tree_add_48_2_groupi_n_418);
 assign csa_tree_add_48_2_groupi_n_803 = ~(csa_tree_add_48_2_groupi_n_728 & csa_tree_add_48_2_groupi_n_419);
 assign csa_tree_add_48_2_groupi_n_802 = ~(csa_tree_add_48_2_groupi_n_728 & csa_tree_add_48_2_groupi_n_448);
 assign csa_tree_add_48_2_groupi_n_801 = ~(csa_tree_add_48_2_groupi_n_730 & csa_tree_add_48_2_groupi_n_467);
 assign csa_tree_add_48_2_groupi_n_800 = ~(csa_tree_add_48_2_groupi_n_730 & csa_tree_add_48_2_groupi_n_474);
 assign csa_tree_add_48_2_groupi_n_799 = ~(csa_tree_add_48_2_groupi_n_721 & csa_tree_add_48_2_groupi_n_452);
 assign csa_tree_add_48_2_groupi_n_798 = ~(csa_tree_add_48_2_groupi_n_728 & csa_tree_add_48_2_groupi_n_482);
 assign csa_tree_add_48_2_groupi_n_797 = ~(csa_tree_add_48_2_groupi_n_724 & csa_tree_add_48_2_groupi_n_492);
 assign csa_tree_add_48_2_groupi_n_796 = ~(csa_tree_add_48_2_groupi_n_125 & ~csa_tree_add_48_2_groupi_n_497);
 assign csa_tree_add_48_2_groupi_n_795 = ~(csa_tree_add_48_2_groupi_n_125 & csa_tree_add_48_2_groupi_n_756);
 assign csa_tree_add_48_2_groupi_n_794 = ~(csa_tree_add_48_2_groupi_n_723 | csa_tree_add_48_2_groupi_n_423);
 assign csa_tree_add_48_2_groupi_n_793 = ~(csa_tree_add_48_2_groupi_n_125 & csa_tree_add_48_2_groupi_n_752);
 assign csa_tree_add_48_2_groupi_n_792 = ~(csa_tree_add_48_2_groupi_n_725 | csa_tree_add_48_2_groupi_n_424);
 assign csa_tree_add_48_2_groupi_n_791 = ~(csa_tree_add_48_2_groupi_n_125 & csa_tree_add_48_2_groupi_n_753);
 assign csa_tree_add_48_2_groupi_n_790 = ~(csa_tree_add_48_2_groupi_n_724 & csa_tree_add_48_2_groupi_n_755);
 assign csa_tree_add_48_2_groupi_n_789 = ~(csa_tree_add_48_2_groupi_n_723 | csa_tree_add_48_2_groupi_n_495);
 assign csa_tree_add_48_2_groupi_n_788 = ~(csa_tree_add_48_2_groupi_n_724 & csa_tree_add_48_2_groupi_n_757);
 assign csa_tree_add_48_2_groupi_n_787 = ~(csa_tree_add_48_2_groupi_n_125 & ~csa_tree_add_48_2_groupi_n_496);
 assign csa_tree_add_48_2_groupi_n_786 = ~(csa_tree_add_48_2_groupi_n_724 & csa_tree_add_48_2_groupi_n_751);
 assign csa_tree_add_48_2_groupi_n_785 = ~(csa_tree_add_48_2_groupi_n_725 | ~csa_tree_add_48_2_groupi_n_493);
 assign csa_tree_add_48_2_groupi_n_784 = ~(csa_tree_add_48_2_groupi_n_724 & csa_tree_add_48_2_groupi_n_759);
 assign csa_tree_add_48_2_groupi_n_783 = ~(csa_tree_add_48_2_groupi_n_724 & ~csa_tree_add_48_2_groupi_n_491);
 assign csa_tree_add_48_2_groupi_n_782 = ~(csa_tree_add_48_2_groupi_n_546 & csa_tree_add_48_2_groupi_n_591);
 assign csa_tree_add_48_2_groupi_n_781 = ~(csa_tree_add_48_2_groupi_n_727 & csa_tree_add_48_2_groupi_n_420);
 assign csa_tree_add_48_2_groupi_n_780 = ~(csa_tree_add_48_2_groupi_n_546 & csa_tree_add_48_2_groupi_n_617);
 assign csa_tree_add_48_2_groupi_n_779 = ~(csa_tree_add_48_2_groupi_n_546 & csa_tree_add_48_2_groupi_n_604);
 assign csa_tree_add_48_2_groupi_n_778 = ~(csa_tree_add_48_2_groupi_n_546 & csa_tree_add_48_2_groupi_n_600);
 assign csa_tree_add_48_2_groupi_n_777 = ~(csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_584);
 assign csa_tree_add_48_2_groupi_n_776 = ~(csa_tree_add_48_2_groupi_n_546 & csa_tree_add_48_2_groupi_n_596);
 assign csa_tree_add_48_2_groupi_n_775 = ~(csa_tree_add_48_2_groupi_n_546 & csa_tree_add_48_2_groupi_n_598);
 assign csa_tree_add_48_2_groupi_n_774 = ~(csa_tree_add_48_2_groupi_n_123 & csa_tree_add_48_2_groupi_n_515);
 assign csa_tree_add_48_2_groupi_n_773 = ~(csa_tree_add_48_2_groupi_n_123 & csa_tree_add_48_2_groupi_n_511);
 assign csa_tree_add_48_2_groupi_n_772 = ~(csa_tree_add_48_2_groupi_n_124 | csa_tree_add_48_2_groupi_n_425);
 assign csa_tree_add_48_2_groupi_n_771 = ~(csa_tree_add_48_2_groupi_n_678 & csa_tree_add_48_2_groupi_n_445);
 assign csa_tree_add_48_2_groupi_n_770 = (csa_tree_add_48_2_groupi_n_121 & csa_tree_add_48_2_groupi_n_443);
 assign csa_tree_add_48_2_groupi_n_769 = ~(csa_tree_add_48_2_groupi_n_121 & csa_tree_add_48_2_groupi_n_441);
 assign csa_tree_add_48_2_groupi_n_768 = ~(csa_tree_add_48_2_groupi_n_121 & csa_tree_add_48_2_groupi_n_623);
 assign csa_tree_add_48_2_groupi_n_767 = ~(csa_tree_add_48_2_groupi_n_121 & csa_tree_add_48_2_groupi_n_620);
 assign csa_tree_add_48_2_groupi_n_766 = ~(csa_tree_add_48_2_groupi_n_122 | csa_tree_add_48_2_groupi_n_426);
 assign csa_tree_add_48_2_groupi_n_765 = ~(csa_tree_add_48_2_groupi_n_681 & csa_tree_add_48_2_groupi_n_617);
 assign csa_tree_add_48_2_groupi_n_764 = ~(csa_tree_add_48_2_groupi_n_681 & csa_tree_add_48_2_groupi_n_428);
 assign csa_tree_add_48_2_groupi_n_763 = ~(csa_tree_add_48_2_groupi_n_681 & csa_tree_add_48_2_groupi_n_600);
 assign csa_tree_add_48_2_groupi_n_762 = ~csa_tree_add_48_2_groupi_n_598;
 assign csa_tree_add_48_2_groupi_n_761 = ~csa_tree_add_48_2_groupi_n_406;
 assign csa_tree_add_48_2_groupi_n_760 = ~csa_tree_add_48_2_groupi_n_604;
 assign csa_tree_add_48_2_groupi_n_758 = ~csa_tree_add_48_2_groupi_n_411;
 assign csa_tree_add_48_2_groupi_n_754 = ~csa_tree_add_48_2_groupi_n_304;
 assign csa_tree_add_48_2_groupi_n_750 = ~csa_tree_add_48_2_groupi_n_405;
 assign csa_tree_add_48_2_groupi_n_749 = ~csa_tree_add_48_2_groupi_n_402;
 assign csa_tree_add_48_2_groupi_n_743 = ~csa_tree_add_48_2_groupi_n_742;
 assign csa_tree_add_48_2_groupi_n_741 = ~csa_tree_add_48_2_groupi_n_740;
 assign csa_tree_add_48_2_groupi_n_739 = ~csa_tree_add_48_2_groupi_n_738;
 assign csa_tree_add_48_2_groupi_n_737 = ~csa_tree_add_48_2_groupi_n_736;
 assign csa_tree_add_48_2_groupi_n_733 = ~csa_tree_add_48_2_groupi_n_732;
 assign csa_tree_add_48_2_groupi_n_729 = ~csa_tree_add_48_2_groupi_n_730;
 assign csa_tree_add_48_2_groupi_n_726 = ~csa_tree_add_48_2_groupi_n_727;
 assign csa_tree_add_48_2_groupi_n_724 = ~csa_tree_add_48_2_groupi_n_725;
 assign csa_tree_add_48_2_groupi_n_723 = ~csa_tree_add_48_2_groupi_n_125;
 assign csa_tree_add_48_2_groupi_n_721 = ~csa_tree_add_48_2_groupi_n_722;
 assign csa_tree_add_48_2_groupi_n_720 = ({in4[7]} & {in3[5]});
 assign csa_tree_add_48_2_groupi_n_759 = ({in4[7]} ^ {in3[5]});
 assign csa_tree_add_48_2_groupi_n_719 = ({in4[7]} & {in3[6]});
 assign csa_tree_add_48_2_groupi_n_757 = ({in4[7]} ^ {in3[6]});
 assign csa_tree_add_48_2_groupi_n_718 = ({in6[7]} & {in5[5]});
 assign csa_tree_add_48_2_groupi_n_756 = ({in6[7]} ^ {in5[5]});
 assign csa_tree_add_48_2_groupi_n_717 = ({in4[7]} & {in3[7]});
 assign csa_tree_add_48_2_groupi_n_755 = ({in4[7]} ^ {in3[7]});
 assign csa_tree_add_48_2_groupi_n_716 = ({in6[7]} & {in5[6]});
 assign csa_tree_add_48_2_groupi_n_753 = ({in6[7]} ^ {in5[6]});
 assign csa_tree_add_48_2_groupi_n_715 = ({in6[7]} & {in5[7]});
 assign csa_tree_add_48_2_groupi_n_752 = ({in6[7]} ^ {in5[7]});
 assign csa_tree_add_48_2_groupi_n_714 = ({in4[7]} & {in3[4]});
 assign csa_tree_add_48_2_groupi_n_751 = ({in4[7]} ^ {in3[4]});
 assign csa_tree_add_48_2_groupi_n_713 = ~(csa_tree_add_48_2_groupi_n_555 | csa_tree_add_48_2_groupi_n_554);
 assign csa_tree_add_48_2_groupi_n_712 = ~(csa_tree_add_48_2_groupi_n_476 | csa_tree_add_48_2_groupi_n_181);
 assign csa_tree_add_48_2_groupi_n_711 = ~(csa_tree_add_48_2_groupi_n_468 & {in6[0]});
 assign csa_tree_add_48_2_groupi_n_748 = ~(csa_tree_add_48_2_groupi_n_458 & {in6[0]});
 assign csa_tree_add_48_2_groupi_n_710 = ~(csa_tree_add_48_2_groupi_n_480 | csa_tree_add_48_2_groupi_n_181);
 assign csa_tree_add_48_2_groupi_n_709 = ~(csa_tree_add_48_2_groupi_n_472 | csa_tree_add_48_2_groupi_n_181);
 assign csa_tree_add_48_2_groupi_n_708 = ~(csa_tree_add_48_2_groupi_n_471 & {in4[0]});
 assign csa_tree_add_48_2_groupi_n_707 = ~(csa_tree_add_48_2_groupi_n_181 | (csa_tree_add_48_2_groupi_n_305
    & csa_tree_add_48_2_groupi_n_306));
 assign csa_tree_add_48_2_groupi_n_706 = ~(csa_tree_add_48_2_groupi_n_486 & ~csa_tree_add_48_2_groupi_n_142);
 assign csa_tree_add_48_2_groupi_n_705 = ~(csa_tree_add_48_2_groupi_n_460 | csa_tree_add_48_2_groupi_n_142);
 assign csa_tree_add_48_2_groupi_n_704 = ~(csa_tree_add_48_2_groupi_n_451 | csa_tree_add_48_2_groupi_n_181);
 assign csa_tree_add_48_2_groupi_n_703 = ~(csa_tree_add_48_2_groupi_n_477 & {in6[0]});
 assign csa_tree_add_48_2_groupi_n_702 = ~(csa_tree_add_48_2_groupi_n_120 & csa_tree_add_48_2_groupi_n_452);
 assign csa_tree_add_48_2_groupi_n_701 = ~(csa_tree_add_48_2_groupi_n_551 & csa_tree_add_48_2_groupi_n_484);
 assign csa_tree_add_48_2_groupi_n_700 = ~(csa_tree_add_48_2_groupi_n_560 & ~csa_tree_add_48_2_groupi_n_172);
 assign csa_tree_add_48_2_groupi_n_699 = ~(csa_tree_add_48_2_groupi_n_579 & {in2[0]});
 assign csa_tree_add_48_2_groupi_n_698 = ~(csa_tree_add_48_2_groupi_n_581 & ~csa_tree_add_48_2_groupi_n_172);
 assign csa_tree_add_48_2_groupi_n_697 = ~(csa_tree_add_48_2_groupi_n_576 | csa_tree_add_48_2_groupi_n_172);
 assign csa_tree_add_48_2_groupi_n_696 = ~(csa_tree_add_48_2_groupi_n_172 | (csa_tree_add_48_2_groupi_n_307
    & csa_tree_add_48_2_groupi_n_415));
 assign csa_tree_add_48_2_groupi_n_695 = ~(csa_tree_add_48_2_groupi_n_570 & ~csa_tree_add_48_2_groupi_n_172);
 assign csa_tree_add_48_2_groupi_n_694 = ~(csa_tree_add_48_2_groupi_n_574 & {in2[0]});
 assign csa_tree_add_48_2_groupi_n_693 = ~(csa_tree_add_48_2_groupi_n_457 | csa_tree_add_48_2_groupi_n_142);
 assign csa_tree_add_48_2_groupi_n_692 = ~(csa_tree_add_48_2_groupi_n_558 | csa_tree_add_48_2_groupi_n_172);
 assign csa_tree_add_48_2_groupi_n_691 = ~(csa_tree_add_48_2_groupi_n_564 & {in2[0]});
 assign csa_tree_add_48_2_groupi_n_690 = ~(csa_tree_add_48_2_groupi_n_582 & {in2[0]});
 assign csa_tree_add_48_2_groupi_n_689 = ~(csa_tree_add_48_2_groupi_n_572 & ~csa_tree_add_48_2_groupi_n_172);
 assign csa_tree_add_48_2_groupi_n_688 = ~(csa_tree_add_48_2_groupi_n_555 & csa_tree_add_48_2_groupi_n_554);
 assign csa_tree_add_48_2_groupi_n_687 = ~(csa_tree_add_48_2_groupi_n_569 & {in2[0]});
 assign csa_tree_add_48_2_groupi_n_686 = ~(csa_tree_add_48_2_groupi_n_562 & {in2[0]});
 assign csa_tree_add_48_2_groupi_n_685 = ~(csa_tree_add_48_2_groupi_n_573 & {in2[0]});
 assign csa_tree_add_48_2_groupi_n_747 = ~(csa_tree_add_48_2_groupi_n_118 | csa_tree_add_48_2_groupi_n_174);
 assign csa_tree_add_48_2_groupi_n_746 = ~(csa_tree_add_48_2_groupi_n_120 & {in6[3]});
 assign csa_tree_add_48_2_groupi_n_745 = ~(csa_tree_add_48_2_groupi_n_547 | csa_tree_add_48_2_groupi_n_141);
 assign csa_tree_add_48_2_groupi_n_744 = ~(csa_tree_add_48_2_groupi_n_551 & ~csa_tree_add_48_2_groupi_n_140);
 assign csa_tree_add_48_2_groupi_n_742 = ~(csa_tree_add_48_2_groupi_n_552 & {in4[7]});
 assign csa_tree_add_48_2_groupi_n_740 = ~(csa_tree_add_48_2_groupi_n_550 & {in6[7]});
 assign csa_tree_add_48_2_groupi_n_738 = ~(csa_tree_add_48_2_groupi_n_118 | csa_tree_add_48_2_groupi_n_178);
 assign csa_tree_add_48_2_groupi_n_684 = ~(csa_tree_add_48_2_groupi_n_551 & {in3[0]});
 assign csa_tree_add_48_2_groupi_n_736 = ~(csa_tree_add_48_2_groupi_n_553 | csa_tree_add_48_2_groupi_n_178);
 assign csa_tree_add_48_2_groupi_n_735 = ~(csa_tree_add_48_2_groupi_n_549 | csa_tree_add_48_2_groupi_n_180);
 assign csa_tree_add_48_2_groupi_n_734 = ~(csa_tree_add_48_2_groupi_n_544 & {in1[0]});
 assign csa_tree_add_48_2_groupi_n_732 = ~(csa_tree_add_48_2_groupi_n_547 | csa_tree_add_48_2_groupi_n_180);
 assign csa_tree_add_48_2_groupi_n_683 = ~(csa_tree_add_48_2_groupi_n_542 & {in1[0]});
 assign csa_tree_add_48_2_groupi_n_731 = ~(csa_tree_add_48_2_groupi_n_545 | csa_tree_add_48_2_groupi_n_179);
 assign csa_tree_add_48_2_groupi_n_682 = ~(csa_tree_add_48_2_groupi_n_120 & {in5[0]});
 assign csa_tree_add_48_2_groupi_n_730 = ~(csa_tree_add_48_2_groupi_n_548 | csa_tree_add_48_2_groupi_n_527);
 assign csa_tree_add_48_2_groupi_n_728 = ~(csa_tree_add_48_2_groupi_n_117 | csa_tree_add_48_2_groupi_n_525);
 assign csa_tree_add_48_2_groupi_n_727 = ~(csa_tree_add_48_2_groupi_n_551 | csa_tree_add_48_2_groupi_n_524);
 assign csa_tree_add_48_2_groupi_n_725 = ~(csa_tree_add_48_2_groupi_n_553 & csa_tree_add_48_2_groupi_n_529);
 assign csa_tree_add_48_2_groupi_n_125 = ~(csa_tree_add_48_2_groupi_n_550 | csa_tree_add_48_2_groupi_n_528);
 assign csa_tree_add_48_2_groupi_n_722 = ~(csa_tree_add_48_2_groupi_n_119 & csa_tree_add_48_2_groupi_n_526);
 assign csa_tree_add_48_2_groupi_n_680 = ~csa_tree_add_48_2_groupi_n_681;
 assign csa_tree_add_48_2_groupi_n_124 = ~csa_tree_add_48_2_groupi_n_123;
 assign csa_tree_add_48_2_groupi_n_679 = ~csa_tree_add_48_2_groupi_n_123;
 assign csa_tree_add_48_2_groupi_n_122 = ~csa_tree_add_48_2_groupi_n_121;
 assign csa_tree_add_48_2_groupi_n_677 = ~(csa_tree_add_48_2_groupi_n_548 & csa_tree_add_48_2_groupi_n_473);
 assign csa_tree_add_48_2_groupi_n_676 = ~(csa_tree_add_48_2_groupi_n_117 & csa_tree_add_48_2_groupi_n_454);
 assign csa_tree_add_48_2_groupi_n_675 = ~(csa_tree_add_48_2_groupi_n_119 | csa_tree_add_48_2_groupi_n_464);
 assign csa_tree_add_48_2_groupi_n_674 = ~(csa_tree_add_48_2_groupi_n_551 & csa_tree_add_48_2_groupi_n_450);
 assign csa_tree_add_48_2_groupi_n_673 = ~(csa_tree_add_48_2_groupi_n_119 | csa_tree_add_48_2_groupi_n_461);
 assign csa_tree_add_48_2_groupi_n_672 = ~(csa_tree_add_48_2_groupi_n_551 & csa_tree_add_48_2_groupi_n_463);
 assign csa_tree_add_48_2_groupi_n_671 = ~(csa_tree_add_48_2_groupi_n_548 & csa_tree_add_48_2_groupi_n_456);
 assign csa_tree_add_48_2_groupi_n_670 = ~(csa_tree_add_48_2_groupi_n_119 | csa_tree_add_48_2_groupi_n_446);
 assign csa_tree_add_48_2_groupi_n_669 = ~(csa_tree_add_48_2_groupi_n_548 & csa_tree_add_48_2_groupi_n_475);
 assign csa_tree_add_48_2_groupi_n_668 = ~(csa_tree_add_48_2_groupi_n_117 & csa_tree_add_48_2_groupi_n_483);
 assign csa_tree_add_48_2_groupi_n_667 = ~(csa_tree_add_48_2_groupi_n_551 & csa_tree_add_48_2_groupi_n_462);
 assign csa_tree_add_48_2_groupi_n_666 = ~(csa_tree_add_48_2_groupi_n_548 & csa_tree_add_48_2_groupi_n_479);
 assign csa_tree_add_48_2_groupi_n_665 = ~(csa_tree_add_48_2_groupi_n_548 & csa_tree_add_48_2_groupi_n_481);
 assign csa_tree_add_48_2_groupi_n_664 = ~(csa_tree_add_48_2_groupi_n_551 & csa_tree_add_48_2_groupi_n_485);
 assign csa_tree_add_48_2_groupi_n_663 = ~(csa_tree_add_48_2_groupi_n_120 & csa_tree_add_48_2_groupi_n_449);
 assign csa_tree_add_48_2_groupi_n_662 = ~(csa_tree_add_48_2_groupi_n_117 & csa_tree_add_48_2_groupi_n_448);
 assign csa_tree_add_48_2_groupi_n_661 = ~(csa_tree_add_48_2_groupi_n_548 & csa_tree_add_48_2_groupi_n_474);
 assign csa_tree_add_48_2_groupi_n_660 = ~(csa_tree_add_48_2_groupi_n_119 | csa_tree_add_48_2_groupi_n_455);
 assign csa_tree_add_48_2_groupi_n_659 = ~(csa_tree_add_48_2_groupi_n_117 & csa_tree_add_48_2_groupi_n_488);
 assign csa_tree_add_48_2_groupi_n_658 = ~(csa_tree_add_48_2_groupi_n_117 & csa_tree_add_48_2_groupi_n_469);
 assign csa_tree_add_48_2_groupi_n_657 = ~(csa_tree_add_48_2_groupi_n_117 & csa_tree_add_48_2_groupi_n_482);
 assign csa_tree_add_48_2_groupi_n_656 = ~(csa_tree_add_48_2_groupi_n_117 & csa_tree_add_48_2_groupi_n_453);
 assign csa_tree_add_48_2_groupi_n_655 = ~(csa_tree_add_48_2_groupi_n_534 & csa_tree_add_48_2_groupi_n_111);
 assign csa_tree_add_48_2_groupi_n_654 = ~(csa_tree_add_48_2_groupi_n_120 & csa_tree_add_48_2_groupi_n_465);
 assign csa_tree_add_48_2_groupi_n_653 = ~(csa_tree_add_48_2_groupi_n_537 | csa_tree_add_48_2_groupi_n_393);
 assign csa_tree_add_48_2_groupi_n_652 = ~(csa_tree_add_48_2_groupi_n_544 & csa_tree_add_48_2_groupi_n_510);
 assign csa_tree_add_48_2_groupi_n_651 = ~(csa_tree_add_48_2_groupi_n_544 & csa_tree_add_48_2_groupi_n_512);
 assign csa_tree_add_48_2_groupi_n_650 = ~(csa_tree_add_48_2_groupi_n_544 & csa_tree_add_48_2_groupi_n_514);
 assign csa_tree_add_48_2_groupi_n_649 = ~(csa_tree_add_48_2_groupi_n_544 & ~csa_tree_add_48_2_groupi_n_498);
 assign csa_tree_add_48_2_groupi_n_648 = ~(csa_tree_add_48_2_groupi_n_544 & csa_tree_add_48_2_groupi_n_515);
 assign csa_tree_add_48_2_groupi_n_647 = ~(csa_tree_add_48_2_groupi_n_543 | csa_tree_add_48_2_groupi_n_518);
 assign csa_tree_add_48_2_groupi_n_646 = ~(csa_tree_add_48_2_groupi_n_544 & csa_tree_add_48_2_groupi_n_505);
 assign csa_tree_add_48_2_groupi_n_645 = ~(csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_624);
 assign csa_tree_add_48_2_groupi_n_644 = ~(csa_tree_add_48_2_groupi_n_542 & csa_tree_add_48_2_groupi_n_630);
 assign csa_tree_add_48_2_groupi_n_643 = ~(csa_tree_add_48_2_groupi_n_542 & csa_tree_add_48_2_groupi_n_445);
 assign csa_tree_add_48_2_groupi_n_642 = ~(csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_605);
 assign csa_tree_add_48_2_groupi_n_641 = ~(csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_444);
 assign csa_tree_add_48_2_groupi_n_640 = ~(csa_tree_add_48_2_groupi_n_542 & csa_tree_add_48_2_groupi_n_623);
 assign csa_tree_add_48_2_groupi_n_639 = ~(csa_tree_add_48_2_groupi_n_542 & csa_tree_add_48_2_groupi_n_620);
 assign csa_tree_add_48_2_groupi_n_638 = ~(csa_tree_add_48_2_groupi_n_542 & csa_tree_add_48_2_groupi_n_434);
 assign csa_tree_add_48_2_groupi_n_637 = ~(csa_tree_add_48_2_groupi_n_541 | ~csa_tree_add_48_2_groupi_n_441);
 assign csa_tree_add_48_2_groupi_n_636 = ~(csa_tree_add_48_2_groupi_n_542 & csa_tree_add_48_2_groupi_n_615);
 assign csa_tree_add_48_2_groupi_n_635 = ~(csa_tree_add_48_2_groupi_n_541 | csa_tree_add_48_2_groupi_n_442);
 assign csa_tree_add_48_2_groupi_n_634 = ~(csa_tree_add_48_2_groupi_n_536 | csa_tree_add_48_2_groupi_n_398);
 assign csa_tree_add_48_2_groupi_n_681 = ~(csa_tree_add_48_2_groupi_n_546 | csa_tree_add_48_2_groupi_n_532);
 assign csa_tree_add_48_2_groupi_n_123 = ~(csa_tree_add_48_2_groupi_n_544 | csa_tree_add_48_2_groupi_n_531);
 assign csa_tree_add_48_2_groupi_n_678 = ~(csa_tree_add_48_2_groupi_n_542 | csa_tree_add_48_2_groupi_n_633);
 assign csa_tree_add_48_2_groupi_n_121 = ~(csa_tree_add_48_2_groupi_n_542 | csa_tree_add_48_2_groupi_n_633);
 assign csa_tree_add_48_2_groupi_n_631 = ~csa_tree_add_48_2_groupi_n_630;
 assign csa_tree_add_48_2_groupi_n_625 = ~csa_tree_add_48_2_groupi_n_624;
 assign csa_tree_add_48_2_groupi_n_616 = ~csa_tree_add_48_2_groupi_n_615;
 assign csa_tree_add_48_2_groupi_n_583 = ~csa_tree_add_48_2_groupi_n_582;
 assign csa_tree_add_48_2_groupi_n_580 = ~csa_tree_add_48_2_groupi_n_579;
 assign csa_tree_add_48_2_groupi_n_575 = ~csa_tree_add_48_2_groupi_n_574;
 assign csa_tree_add_48_2_groupi_n_565 = ~csa_tree_add_48_2_groupi_n_564;
 assign csa_tree_add_48_2_groupi_n_561 = ~csa_tree_add_48_2_groupi_n_560;
 assign csa_tree_add_48_2_groupi_n_120 = ~csa_tree_add_48_2_groupi_n_119;
 assign csa_tree_add_48_2_groupi_n_552 = ~csa_tree_add_48_2_groupi_n_553;
 assign csa_tree_add_48_2_groupi_n_549 = ~csa_tree_add_48_2_groupi_n_550;
 assign csa_tree_add_48_2_groupi_n_548 = ~csa_tree_add_48_2_groupi_n_118;
 assign csa_tree_add_48_2_groupi_n_545 = ~csa_tree_add_48_2_groupi_n_546;
 assign csa_tree_add_48_2_groupi_n_543 = ~csa_tree_add_48_2_groupi_n_544;
 assign csa_tree_add_48_2_groupi_n_541 = ~csa_tree_add_48_2_groupi_n_542;
 assign csa_tree_add_48_2_groupi_n_540 = ~(csa_tree_add_48_2_groupi_n_396 & csa_tree_add_48_2_groupi_n_174);
 assign csa_tree_add_48_2_groupi_n_539 = ~(csa_tree_add_48_2_groupi_n_401 & csa_tree_add_48_2_groupi_n_141);
 assign csa_tree_add_48_2_groupi_n_538 = ~({in4[3]} | ({in4[4]} & {in3[0]}));
 assign csa_tree_add_48_2_groupi_n_537 = ~({in6[1]} | ({in6[2]} & {in5[0]}));
 assign csa_tree_add_48_2_groupi_n_536 = ~({in4[1]} | ({in4[2]} & {in3[0]}));
 assign csa_tree_add_48_2_groupi_n_535 = ~(csa_tree_add_48_2_groupi_n_394 & csa_tree_add_48_2_groupi_n_138);
 assign csa_tree_add_48_2_groupi_n_534 = ~(csa_tree_add_48_2_groupi_n_397 & csa_tree_add_48_2_groupi_n_171);
 assign csa_tree_add_48_2_groupi_n_533 = ~({in2[1]} | ({in2[2]} & {in1[0]}));
 assign csa_tree_add_48_2_groupi_n_532 = ~(csa_tree_add_48_2_groupi_n_362 | csa_tree_add_48_2_groupi_n_354);
 assign csa_tree_add_48_2_groupi_n_633 = ~(csa_tree_add_48_2_groupi_n_348 | csa_tree_add_48_2_groupi_n_351);
 assign csa_tree_add_48_2_groupi_n_531 = ~(csa_tree_add_48_2_groupi_n_370 | csa_tree_add_48_2_groupi_n_383);
 assign csa_tree_add_48_2_groupi_n_530 = ~({in2[5]} ^ {in1[27]});
 assign csa_tree_add_48_2_groupi_n_529 = ~(csa_tree_add_48_2_groupi_n_361 & csa_tree_add_48_2_groupi_n_349);
 assign csa_tree_add_48_2_groupi_n_528 = ~(csa_tree_add_48_2_groupi_n_358 | csa_tree_add_48_2_groupi_n_380);
 assign csa_tree_add_48_2_groupi_n_527 = ~(csa_tree_add_48_2_groupi_n_353 | csa_tree_add_48_2_groupi_n_364);
 assign csa_tree_add_48_2_groupi_n_526 = ~(csa_tree_add_48_2_groupi_n_356 & csa_tree_add_48_2_groupi_n_372);
 assign csa_tree_add_48_2_groupi_n_525 = ~(csa_tree_add_48_2_groupi_n_359 | csa_tree_add_48_2_groupi_n_379);
 assign csa_tree_add_48_2_groupi_n_524 = ~(csa_tree_add_48_2_groupi_n_355 | csa_tree_add_48_2_groupi_n_350);
 assign csa_tree_add_48_2_groupi_n_523 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[25]}) | (csa_tree_add_48_2_groupi_n_197
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_522 = ~({in6[3]} | ({in6[4]} & {in5[0]}));
 assign csa_tree_add_48_2_groupi_n_632 = ~({in2[5]} ^ {in1[26]});
 assign csa_tree_add_48_2_groupi_n_630 = ~((csa_tree_add_48_2_groupi_n_186 & ~{in2[3]}) | ({in1[12]}
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_629 = ~({in2[1]} ^ {in1[26]});
 assign csa_tree_add_48_2_groupi_n_628 = ~({in2[1]} ^ {in1[28]});
 assign csa_tree_add_48_2_groupi_n_627 = ~({in2[1]} ^ {in1[27]});
 assign csa_tree_add_48_2_groupi_n_626 = ~((csa_tree_add_48_2_groupi_n_171 & {in1[13]}) | (csa_tree_add_48_2_groupi_n_195
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_624 = ~(({in1[8]} & ~{in2[3]}) | (csa_tree_add_48_2_groupi_n_143 &
    {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_623 = ~(csa_tree_add_48_2_groupi_n_243 & ~(csa_tree_add_48_2_groupi_n_171
    & {in1[9]}));
 assign csa_tree_add_48_2_groupi_n_622 = ~(({in2[3]} & ~{in1[28]}) | (csa_tree_add_48_2_groupi_n_171
    & {in1[28]}));
 assign csa_tree_add_48_2_groupi_n_621 = ~((csa_tree_add_48_2_groupi_n_171 & {in1[23]}) | (csa_tree_add_48_2_groupi_n_153
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_620 = ~((csa_tree_add_48_2_groupi_n_189 & ~{in2[3]}) | ({in1[6]} &
    {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_619 = ~((csa_tree_add_48_2_groupi_n_171 & {in1[20]}) | (csa_tree_add_48_2_groupi_n_193
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_618 = ~(({in2[3]} & ~{in1[27]}) | (csa_tree_add_48_2_groupi_n_171
    & {in1[27]}));
 assign csa_tree_add_48_2_groupi_n_617 = ~(csa_tree_add_48_2_groupi_n_266 & csa_tree_add_48_2_groupi_n_273);
 assign csa_tree_add_48_2_groupi_n_615 = ~(csa_tree_add_48_2_groupi_n_223 & csa_tree_add_48_2_groupi_n_268);
 assign csa_tree_add_48_2_groupi_n_614 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[24]}) | (csa_tree_add_48_2_groupi_n_165
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_613 = ~(({in2[3]} & ~{in1[26]}) | (csa_tree_add_48_2_groupi_n_171
    & {in1[26]}));
 assign csa_tree_add_48_2_groupi_n_612 = ~((csa_tree_add_48_2_groupi_n_137 & {in1[25]}) | (csa_tree_add_48_2_groupi_n_197
    & {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_611 = ~((csa_tree_add_48_2_groupi_n_137 & {in1[24]}) | (csa_tree_add_48_2_groupi_n_165
    & {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_610 = ~((csa_tree_add_48_2_groupi_n_171 & {in1[24]}) | (csa_tree_add_48_2_groupi_n_165
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_609 = ~((csa_tree_add_48_2_groupi_n_171 & {in1[25]}) | (csa_tree_add_48_2_groupi_n_197
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_608 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[24]}) | (csa_tree_add_48_2_groupi_n_165
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_607 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[25]}) | (csa_tree_add_48_2_groupi_n_197
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_606 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[22]}) | (csa_tree_add_48_2_groupi_n_145
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_605 = ~(({in1[4]} & ~{in2[3]}) | (csa_tree_add_48_2_groupi_n_157 &
    {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_604 = ~((csa_tree_add_48_2_groupi_n_143 & ~{in2[7]}) | ({in1[8]} &
    {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_603 = ~((csa_tree_add_48_2_groupi_n_149 & ~{in2[7]}) | ({in1[5]} &
    {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_602 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[10]}) | (csa_tree_add_48_2_groupi_n_185
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_601 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[23]}) | (csa_tree_add_48_2_groupi_n_153
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_600 = ~(csa_tree_add_48_2_groupi_n_263 & csa_tree_add_48_2_groupi_n_289);
 assign csa_tree_add_48_2_groupi_n_599 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[21]}) | (csa_tree_add_48_2_groupi_n_160
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_598 = ~(csa_tree_add_48_2_groupi_n_385 & csa_tree_add_48_2_groupi_n_242);
 assign csa_tree_add_48_2_groupi_n_597 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[15]}) | (csa_tree_add_48_2_groupi_n_156
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_596 = ~((csa_tree_add_48_2_groupi_n_182 & ~{in2[7]}) | ({in1[7]} &
    {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_595 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[13]}) | (csa_tree_add_48_2_groupi_n_195
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_594 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[16]}) | (csa_tree_add_48_2_groupi_n_152
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_593 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[19]}) | (csa_tree_add_48_2_groupi_n_159
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_592 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[18]}) | (csa_tree_add_48_2_groupi_n_150
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_591 = ~((csa_tree_add_48_2_groupi_n_189 & ~{in2[7]}) | ({in1[6]} &
    {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_590 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[9]}) | (csa_tree_add_48_2_groupi_n_148
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_589 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[11]}) | (csa_tree_add_48_2_groupi_n_196
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_588 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[17]}) | (csa_tree_add_48_2_groupi_n_154
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_587 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[12]}) | (csa_tree_add_48_2_groupi_n_186
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_586 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[20]}) | (csa_tree_add_48_2_groupi_n_193
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_585 = ~((csa_tree_add_48_2_groupi_n_136 & {in1[14]}) | (csa_tree_add_48_2_groupi_n_164
    & {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_584 = ~(({in1[4]} & ~{in2[7]}) | (csa_tree_add_48_2_groupi_n_157 &
    {in2[7]}));
 assign csa_tree_add_48_2_groupi_n_582 = ~(csa_tree_add_48_2_groupi_n_221 & csa_tree_add_48_2_groupi_n_389);
 assign csa_tree_add_48_2_groupi_n_581 = ~((csa_tree_add_48_2_groupi_n_182 & ~{in2[1]}) | ({in1[7]} &
    {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_579 = ~(csa_tree_add_48_2_groupi_n_271 & ~(csa_tree_add_48_2_groupi_n_137
    & {in1[14]}));
 assign csa_tree_add_48_2_groupi_n_578 = ~((csa_tree_add_48_2_groupi_n_137 & {in1[23]}) | (csa_tree_add_48_2_groupi_n_153
    & {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_577 = ~((csa_tree_add_48_2_groupi_n_137 & {in1[22]}) | (csa_tree_add_48_2_groupi_n_145
    & {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_576 = ~(({in1[6]} & ~{in2[1]}) | (csa_tree_add_48_2_groupi_n_189 &
    {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_574 = ~(csa_tree_add_48_2_groupi_n_276 & csa_tree_add_48_2_groupi_n_345);
 assign csa_tree_add_48_2_groupi_n_573 = ~(({in2[1]} | csa_tree_add_48_2_groupi_n_143) & ({in1[8]} |
    csa_tree_add_48_2_groupi_n_137));
 assign csa_tree_add_48_2_groupi_n_572 = ~((csa_tree_add_48_2_groupi_n_195 & ~{in2[1]}) | ({in1[13]}
    & {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_571 = ~((csa_tree_add_48_2_groupi_n_137 & {in1[16]}) | (csa_tree_add_48_2_groupi_n_152
    & {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_570 = ~((csa_tree_add_48_2_groupi_n_186 & ~{in2[1]}) | ({in1[12]}
    & {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_569 = ~(csa_tree_add_48_2_groupi_n_258 & csa_tree_add_48_2_groupi_n_301);
 assign csa_tree_add_48_2_groupi_n_521 = ~(csa_tree_add_48_2_groupi_n_307 & csa_tree_add_48_2_groupi_n_415);
 assign csa_tree_add_48_2_groupi_n_568 = ~((csa_tree_add_48_2_groupi_n_137 & {in1[20]}) | (csa_tree_add_48_2_groupi_n_193
    & {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_567 = ~((csa_tree_add_48_2_groupi_n_137 & {in1[21]}) | (csa_tree_add_48_2_groupi_n_160
    & {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_566 = ~((csa_tree_add_48_2_groupi_n_137 & {in1[18]}) | (csa_tree_add_48_2_groupi_n_150
    & {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_564 = ~(csa_tree_add_48_2_groupi_n_255 & csa_tree_add_48_2_groupi_n_281);
 assign csa_tree_add_48_2_groupi_n_563 = ~((csa_tree_add_48_2_groupi_n_137 & {in1[19]}) | (csa_tree_add_48_2_groupi_n_159
    & {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_562 = ~(csa_tree_add_48_2_groupi_n_224 & csa_tree_add_48_2_groupi_n_293);
 assign csa_tree_add_48_2_groupi_n_560 = ~(csa_tree_add_48_2_groupi_n_299 & csa_tree_add_48_2_groupi_n_303);
 assign csa_tree_add_48_2_groupi_n_559 = ~((csa_tree_add_48_2_groupi_n_137 & {in1[15]}) | (csa_tree_add_48_2_groupi_n_156
    & {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_558 = ~(csa_tree_add_48_2_groupi_n_300 | csa_tree_add_48_2_groupi_n_265);
 assign csa_tree_add_48_2_groupi_n_557 = ~((csa_tree_add_48_2_groupi_n_137 & {in1[17]}) | (csa_tree_add_48_2_groupi_n_154
    & {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_556 = ~(csa_tree_add_48_2_groupi_n_109 | csa_tree_add_48_2_groupi_n_137);
 assign csa_tree_add_48_2_groupi_n_555 = ~(csa_tree_add_48_2_groupi_n_407 & {in4[1]});
 assign csa_tree_add_48_2_groupi_n_554 = ~(csa_tree_add_48_2_groupi_n_403 & {in6[1]});
 assign csa_tree_add_48_2_groupi_n_119 = ~(csa_tree_add_48_2_groupi_n_368 | csa_tree_add_48_2_groupi_n_369);
 assign csa_tree_add_48_2_groupi_n_553 = ~(csa_tree_add_48_2_groupi_n_360 | csa_tree_add_48_2_groupi_n_371);
 assign csa_tree_add_48_2_groupi_n_551 = ~(csa_tree_add_48_2_groupi_n_381 & csa_tree_add_48_2_groupi_n_373);
 assign csa_tree_add_48_2_groupi_n_550 = ~(csa_tree_add_48_2_groupi_n_377 & csa_tree_add_48_2_groupi_n_375);
 assign csa_tree_add_48_2_groupi_n_118 = ~(csa_tree_add_48_2_groupi_n_352 | csa_tree_add_48_2_groupi_n_365);
 assign csa_tree_add_48_2_groupi_n_547 = ~(csa_tree_add_48_2_groupi_n_346 | csa_tree_add_48_2_groupi_n_367);
 assign csa_tree_add_48_2_groupi_n_117 = ~(csa_tree_add_48_2_groupi_n_347 & csa_tree_add_48_2_groupi_n_366);
 assign csa_tree_add_48_2_groupi_n_546 = ~(csa_tree_add_48_2_groupi_n_382 & csa_tree_add_48_2_groupi_n_357);
 assign csa_tree_add_48_2_groupi_n_544 = ~(csa_tree_add_48_2_groupi_n_376 & csa_tree_add_48_2_groupi_n_374);
 assign csa_tree_add_48_2_groupi_n_542 = ~(csa_tree_add_48_2_groupi_n_363 & csa_tree_add_48_2_groupi_n_378);
 assign csa_tree_add_48_2_groupi_n_487 = ~csa_tree_add_48_2_groupi_n_486;
 assign csa_tree_add_48_2_groupi_n_478 = ~csa_tree_add_48_2_groupi_n_477;
 assign csa_tree_add_48_2_groupi_n_459 = ~csa_tree_add_48_2_groupi_n_458;
 assign csa_tree_add_48_2_groupi_n_447 = ~csa_tree_add_48_2_groupi_n_446;
 assign csa_tree_add_48_2_groupi_n_430 = ~(({in3[0]} & ~{in4[1]}) | (csa_tree_add_48_2_groupi_n_178 &
    {in4[1]}));
 assign csa_tree_add_48_2_groupi_n_428 = ~(csa_tree_add_48_2_groupi_n_203 & csa_tree_add_48_2_groupi_n_204);
 assign csa_tree_add_48_2_groupi_n_427 = ~(({in1[0]} & ~{in2[1]}) | (csa_tree_add_48_2_groupi_n_179 &
    {in2[1]}));
 assign csa_tree_add_48_2_groupi_n_426 = ~(({in1[0]} & ~{in2[3]}) | (csa_tree_add_48_2_groupi_n_179 &
    {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_425 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[0]}) | (csa_tree_add_48_2_groupi_n_179
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_424 = ~(({in4[7]} & ~{in3[0]}) | (csa_tree_add_48_2_groupi_n_173 &
    {in3[0]}));
 assign csa_tree_add_48_2_groupi_n_423 = ~(csa_tree_add_48_2_groupi_n_210 | csa_tree_add_48_2_groupi_n_216);
 assign csa_tree_add_48_2_groupi_n_422 = ~(({in5[0]} & ~{in6[1]}) | (csa_tree_add_48_2_groupi_n_180 &
    {in6[1]}));
 assign csa_tree_add_48_2_groupi_n_421 = ~(csa_tree_add_48_2_groupi_n_207 & csa_tree_add_48_2_groupi_n_211);
 assign csa_tree_add_48_2_groupi_n_420 = ~(csa_tree_add_48_2_groupi_n_208 & csa_tree_add_48_2_groupi_n_209);
 assign csa_tree_add_48_2_groupi_n_419 = ~(csa_tree_add_48_2_groupi_n_206 & csa_tree_add_48_2_groupi_n_205);
 assign csa_tree_add_48_2_groupi_n_418 = ~((csa_tree_add_48_2_groupi_n_174 & ~{in3[0]}) | ({in4[5]} &
    {in3[0]}));
 assign csa_tree_add_48_2_groupi_n_520 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[22]}) | (csa_tree_add_48_2_groupi_n_145
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_519 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[16]}) | (csa_tree_add_48_2_groupi_n_152
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_518 = ~(({in1[3]} & ~{in2[5]}) | (csa_tree_add_48_2_groupi_n_163 &
    {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_517 = ~((csa_tree_add_48_2_groupi_n_182 & ~{in2[5]}) | ({in1[7]} &
    {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_516 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[11]}) | (csa_tree_add_48_2_groupi_n_196
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_515 = ~((csa_tree_add_48_2_groupi_n_157 & ~{in2[5]}) | ({in1[4]} &
    {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_514 = ~((csa_tree_add_48_2_groupi_n_189 & ~{in2[5]}) | ({in1[6]} &
    {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_513 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[17]}) | (csa_tree_add_48_2_groupi_n_154
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_512 = ~((csa_tree_add_48_2_groupi_n_143 & ~{in2[5]}) | ({in1[8]} &
    {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_511 = ~(csa_tree_add_48_2_groupi_n_239 & csa_tree_add_48_2_groupi_n_298);
 assign csa_tree_add_48_2_groupi_n_510 = ~(csa_tree_add_48_2_groupi_n_246 & csa_tree_add_48_2_groupi_n_222);
 assign csa_tree_add_48_2_groupi_n_509 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[18]}) | (csa_tree_add_48_2_groupi_n_150
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_508 = ~(({in1[2]} & ~{in2[5]}) | (csa_tree_add_48_2_groupi_n_158 &
    {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_507 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[21]}) | (csa_tree_add_48_2_groupi_n_160
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_506 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[23]}) | (csa_tree_add_48_2_groupi_n_153
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_505 = ~((csa_tree_add_48_2_groupi_n_148 & ~{in2[5]}) | ({in1[9]} &
    {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_504 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[19]}) | (csa_tree_add_48_2_groupi_n_159
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_503 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[14]}) | (csa_tree_add_48_2_groupi_n_164
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_502 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[20]}) | (csa_tree_add_48_2_groupi_n_193
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_501 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[13]}) | (csa_tree_add_48_2_groupi_n_195
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_500 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[12]}) | (csa_tree_add_48_2_groupi_n_186
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_499 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[15]}) | (csa_tree_add_48_2_groupi_n_156
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_498 = ~((csa_tree_add_48_2_groupi_n_138 & {in1[10]}) | (csa_tree_add_48_2_groupi_n_185
    & {in2[5]}));
 assign csa_tree_add_48_2_groupi_n_497 = ~(csa_tree_add_48_2_groupi_n_252 | csa_tree_add_48_2_groupi_n_332);
 assign csa_tree_add_48_2_groupi_n_496 = ~(({in5[4]} & ~{in6[7]}) | (csa_tree_add_48_2_groupi_n_155 &
    {in6[7]}));
 assign csa_tree_add_48_2_groupi_n_495 = ~((csa_tree_add_48_2_groupi_n_139 & {in5[3]}) | (csa_tree_add_48_2_groupi_n_192
    & {in6[7]}));
 assign csa_tree_add_48_2_groupi_n_494 = ~(csa_tree_add_48_2_groupi_n_392 & csa_tree_add_48_2_groupi_n_251);
 assign csa_tree_add_48_2_groupi_n_493 = ~(csa_tree_add_48_2_groupi_n_285 & csa_tree_add_48_2_groupi_n_245);
 assign csa_tree_add_48_2_groupi_n_492 = ~(csa_tree_add_48_2_groupi_n_339 & csa_tree_add_48_2_groupi_n_235);
 assign csa_tree_add_48_2_groupi_n_491 = ~(({in3[1]} & ~{in4[7]}) | (csa_tree_add_48_2_groupi_n_162 &
    {in4[7]}));
 assign csa_tree_add_48_2_groupi_n_490 = ~(csa_tree_add_48_2_groupi_n_390 | csa_tree_add_48_2_groupi_n_277);
 assign csa_tree_add_48_2_groupi_n_489 = ~(({in3[7]} & ~{in4[1]}) | (csa_tree_add_48_2_groupi_n_187 &
    {in4[1]}));
 assign csa_tree_add_48_2_groupi_n_488 = ~(csa_tree_add_48_2_groupi_n_260 & csa_tree_add_48_2_groupi_n_247);
 assign csa_tree_add_48_2_groupi_n_486 = ~(csa_tree_add_48_2_groupi_n_342 & csa_tree_add_48_2_groupi_n_264);
 assign csa_tree_add_48_2_groupi_n_485 = ~(csa_tree_add_48_2_groupi_n_254 & csa_tree_add_48_2_groupi_n_220);
 assign csa_tree_add_48_2_groupi_n_484 = ~(csa_tree_add_48_2_groupi_n_286 & csa_tree_add_48_2_groupi_n_230);
 assign csa_tree_add_48_2_groupi_n_483 = ~(csa_tree_add_48_2_groupi_n_237 & csa_tree_add_48_2_groupi_n_232);
 assign csa_tree_add_48_2_groupi_n_482 = ~(csa_tree_add_48_2_groupi_n_337 & csa_tree_add_48_2_groupi_n_333);
 assign csa_tree_add_48_2_groupi_n_481 = ~(csa_tree_add_48_2_groupi_n_344 & csa_tree_add_48_2_groupi_n_335);
 assign csa_tree_add_48_2_groupi_n_480 = ~(csa_tree_add_48_2_groupi_n_249 | csa_tree_add_48_2_groupi_n_219);
 assign csa_tree_add_48_2_groupi_n_479 = ~(csa_tree_add_48_2_groupi_n_233 & csa_tree_add_48_2_groupi_n_338);
 assign csa_tree_add_48_2_groupi_n_416 = ~(csa_tree_add_48_2_groupi_n_305 & csa_tree_add_48_2_groupi_n_306);
 assign csa_tree_add_48_2_groupi_n_477 = ~(csa_tree_add_48_2_groupi_n_228 & csa_tree_add_48_2_groupi_n_282);
 assign csa_tree_add_48_2_groupi_n_476 = ~(csa_tree_add_48_2_groupi_n_388 | csa_tree_add_48_2_groupi_n_226);
 assign csa_tree_add_48_2_groupi_n_475 = ~(csa_tree_add_48_2_groupi_n_240 & csa_tree_add_48_2_groupi_n_238);
 assign csa_tree_add_48_2_groupi_n_474 = ~(csa_tree_add_48_2_groupi_n_261 & csa_tree_add_48_2_groupi_n_272);
 assign csa_tree_add_48_2_groupi_n_473 = ~(csa_tree_add_48_2_groupi_n_279 & csa_tree_add_48_2_groupi_n_262);
 assign csa_tree_add_48_2_groupi_n_472 = ~(csa_tree_add_48_2_groupi_n_294 | csa_tree_add_48_2_groupi_n_270);
 assign csa_tree_add_48_2_groupi_n_471 = ~(csa_tree_add_48_2_groupi_n_274 & csa_tree_add_48_2_groupi_n_288);
 assign csa_tree_add_48_2_groupi_n_470 = ~(({in3[3]} & ~{in4[3]}) | (csa_tree_add_48_2_groupi_n_191 &
    {in4[3]}));
 assign csa_tree_add_48_2_groupi_n_469 = ~(csa_tree_add_48_2_groupi_n_340 & csa_tree_add_48_2_groupi_n_227);
 assign csa_tree_add_48_2_groupi_n_468 = ~(csa_tree_add_48_2_groupi_n_296 & csa_tree_add_48_2_groupi_n_384);
 assign csa_tree_add_48_2_groupi_n_467 = ~(csa_tree_add_48_2_groupi_n_391 & csa_tree_add_48_2_groupi_n_250);
 assign csa_tree_add_48_2_groupi_n_466 = ~(({in3[2]} & ~{in4[3]}) | (csa_tree_add_48_2_groupi_n_184 &
    {in4[3]}));
 assign csa_tree_add_48_2_groupi_n_465 = ~(csa_tree_add_48_2_groupi_n_225 & csa_tree_add_48_2_groupi_n_334);
 assign csa_tree_add_48_2_groupi_n_464 = ~(({in5[3]} & ~{in6[3]}) | (csa_tree_add_48_2_groupi_n_192 &
    {in6[3]}));
 assign csa_tree_add_48_2_groupi_n_463 = ~(csa_tree_add_48_2_groupi_n_336 & csa_tree_add_48_2_groupi_n_341);
 assign csa_tree_add_48_2_groupi_n_462 = ~(csa_tree_add_48_2_groupi_n_234 & csa_tree_add_48_2_groupi_n_290);
 assign csa_tree_add_48_2_groupi_n_461 = ~(({in5[2]} & ~{in6[3]}) | (csa_tree_add_48_2_groupi_n_144 &
    {in6[3]}));
 assign csa_tree_add_48_2_groupi_n_460 = ~(csa_tree_add_48_2_groupi_n_295 | csa_tree_add_48_2_groupi_n_287);
 assign csa_tree_add_48_2_groupi_n_458 = ~(csa_tree_add_48_2_groupi_n_291 & csa_tree_add_48_2_groupi_n_280);
 assign csa_tree_add_48_2_groupi_n_457 = ~(csa_tree_add_48_2_groupi_n_275 | csa_tree_add_48_2_groupi_n_283);
 assign csa_tree_add_48_2_groupi_n_456 = ~(csa_tree_add_48_2_groupi_n_244 & csa_tree_add_48_2_groupi_n_229);
 assign csa_tree_add_48_2_groupi_n_455 = ~(csa_tree_add_48_2_groupi_n_248 | csa_tree_add_48_2_groupi_n_253);
 assign csa_tree_add_48_2_groupi_n_454 = ~(csa_tree_add_48_2_groupi_n_278 & csa_tree_add_48_2_groupi_n_267);
 assign csa_tree_add_48_2_groupi_n_453 = ~(csa_tree_add_48_2_groupi_n_331 & csa_tree_add_48_2_groupi_n_269);
 assign csa_tree_add_48_2_groupi_n_452 = ~(csa_tree_add_48_2_groupi_n_257 & ~(csa_tree_add_48_2_groupi_n_175
    & {in5[7]}));
 assign csa_tree_add_48_2_groupi_n_451 = ~(csa_tree_add_48_2_groupi_n_236 | csa_tree_add_48_2_groupi_n_259);
 assign csa_tree_add_48_2_groupi_n_450 = ~(csa_tree_add_48_2_groupi_n_386 & csa_tree_add_48_2_groupi_n_284);
 assign csa_tree_add_48_2_groupi_n_449 = ~(csa_tree_add_48_2_groupi_n_343 & csa_tree_add_48_2_groupi_n_387);
 assign csa_tree_add_48_2_groupi_n_448 = ~(csa_tree_add_48_2_groupi_n_297 & csa_tree_add_48_2_groupi_n_241);
 assign csa_tree_add_48_2_groupi_n_446 = ~(csa_tree_add_48_2_groupi_n_256 | csa_tree_add_48_2_groupi_n_302);
 assign csa_tree_add_48_2_groupi_n_445 = ~((csa_tree_add_48_2_groupi_n_149 & ~{in2[3]}) | ({in1[5]} &
    {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_444 = ~((csa_tree_add_48_2_groupi_n_171 & {in1[3]}) | (csa_tree_add_48_2_groupi_n_163
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_443 = ~(csa_tree_add_48_2_groupi_n_231 & csa_tree_add_48_2_groupi_n_292);
 assign csa_tree_add_48_2_groupi_n_442 = ~(({in1[1]} & ~{in2[3]}) | (csa_tree_add_48_2_groupi_n_194 &
    {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_441 = ~((csa_tree_add_48_2_groupi_n_196 & ~{in2[3]}) | ({in1[11]}
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_440 = ~((csa_tree_add_48_2_groupi_n_171 & {in1[15]}) | (csa_tree_add_48_2_groupi_n_156
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_439 = ~((csa_tree_add_48_2_groupi_n_171 & {in1[19]}) | (csa_tree_add_48_2_groupi_n_159
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_438 = ~((csa_tree_add_48_2_groupi_n_171 & {in1[18]}) | (csa_tree_add_48_2_groupi_n_150
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_436 = ~((csa_tree_add_48_2_groupi_n_171 & {in1[21]}) | (csa_tree_add_48_2_groupi_n_160
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_435 = ~((csa_tree_add_48_2_groupi_n_171 & {in1[16]}) | (csa_tree_add_48_2_groupi_n_152
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_434 = ~((csa_tree_add_48_2_groupi_n_185 & ~{in2[3]}) | ({in1[10]}
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_433 = ~((csa_tree_add_48_2_groupi_n_171 & {in1[22]}) | (csa_tree_add_48_2_groupi_n_145
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_432 = ~((csa_tree_add_48_2_groupi_n_171 & {in1[17]}) | (csa_tree_add_48_2_groupi_n_154
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_431 = ~((csa_tree_add_48_2_groupi_n_171 & {in1[14]}) | (csa_tree_add_48_2_groupi_n_164
    & {in2[3]}));
 assign csa_tree_add_48_2_groupi_n_408 = ~csa_tree_add_48_2_groupi_n_407;
 assign csa_tree_add_48_2_groupi_n_404 = ~csa_tree_add_48_2_groupi_n_403;
 assign csa_tree_add_48_2_groupi_n_401 = ~({in6[6]} & {in5[0]});
 assign csa_tree_add_48_2_groupi_n_400 = ~({in4[4]} | {in3[0]});
 assign csa_tree_add_48_2_groupi_n_399 = ~({in6[4]} | {in5[0]});
 assign csa_tree_add_48_2_groupi_n_398 = ~({in4[2]} | {in3[0]});
 assign csa_tree_add_48_2_groupi_n_397 = ~({in2[4]} & {in1[0]});
 assign csa_tree_add_48_2_groupi_n_396 = ~({in4[6]} & {in3[0]});
 assign csa_tree_add_48_2_groupi_n_395 = ~({in2[2]} | {in1[0]});
 assign csa_tree_add_48_2_groupi_n_394 = ~({in2[6]} & {in1[0]});
 assign csa_tree_add_48_2_groupi_n_393 = ~({in6[2]} | {in5[0]});
 assign csa_tree_add_48_2_groupi_n_392 = ~(csa_tree_add_48_2_groupi_n_139 & {in5[2]});
 assign csa_tree_add_48_2_groupi_n_391 = ~(csa_tree_add_48_2_groupi_n_174 & {in3[5]});
 assign csa_tree_add_48_2_groupi_n_390 = ~({in6[1]} | csa_tree_add_48_2_groupi_n_144);
 assign csa_tree_add_48_2_groupi_n_389 = ~(csa_tree_add_48_2_groupi_n_194 & {in2[1]});
 assign csa_tree_add_48_2_groupi_n_388 = ~({in4[1]} | csa_tree_add_48_2_groupi_n_162);
 assign csa_tree_add_48_2_groupi_n_387 = ~(csa_tree_add_48_2_groupi_n_147 & {in6[3]});
 assign csa_tree_add_48_2_groupi_n_386 = ~(csa_tree_add_48_2_groupi_n_140 & {in3[7]});
 assign csa_tree_add_48_2_groupi_n_385 = ~(csa_tree_add_48_2_groupi_n_136 & {in1[3]});
 assign csa_tree_add_48_2_groupi_n_384 = ~(csa_tree_add_48_2_groupi_n_155 & {in6[1]});
 assign csa_tree_add_48_2_groupi_n_383 = ~({in2[5]} | csa_tree_add_48_2_groupi_n_169);
 assign csa_tree_add_48_2_groupi_n_382 = ~(csa_tree_add_48_2_groupi_n_138 & {in2[6]});
 assign csa_tree_add_48_2_groupi_n_381 = ~(csa_tree_add_48_2_groupi_n_176 & {in4[2]});
 assign csa_tree_add_48_2_groupi_n_380 = ~({in6[7]} | csa_tree_add_48_2_groupi_n_200);
 assign csa_tree_add_48_2_groupi_n_379 = ~({in6[5]} | csa_tree_add_48_2_groupi_n_170);
 assign csa_tree_add_48_2_groupi_n_378 = ~(csa_tree_add_48_2_groupi_n_198 & {in2[1]});
 assign csa_tree_add_48_2_groupi_n_377 = ~(csa_tree_add_48_2_groupi_n_141 & {in6[6]});
 assign csa_tree_add_48_2_groupi_n_376 = ~(csa_tree_add_48_2_groupi_n_171 & {in2[4]});
 assign csa_tree_add_48_2_groupi_n_375 = ~(csa_tree_add_48_2_groupi_n_200 & {in6[5]});
 assign csa_tree_add_48_2_groupi_n_374 = ~(csa_tree_add_48_2_groupi_n_169 & {in2[3]});
 assign csa_tree_add_48_2_groupi_n_373 = ~(csa_tree_add_48_2_groupi_n_199 & {in4[1]});
 assign csa_tree_add_48_2_groupi_n_372 = ~(csa_tree_add_48_2_groupi_n_175 & {in6[2]});
 assign csa_tree_add_48_2_groupi_n_371 = ~({in4[6]} | csa_tree_add_48_2_groupi_n_174);
 assign csa_tree_add_48_2_groupi_n_370 = ~({in2[4]} | csa_tree_add_48_2_groupi_n_138);
 assign csa_tree_add_48_2_groupi_n_369 = ~({in6[2]} | csa_tree_add_48_2_groupi_n_177);
 assign csa_tree_add_48_2_groupi_n_368 = ~({in6[1]} | csa_tree_add_48_2_groupi_n_201);
 assign csa_tree_add_48_2_groupi_n_367 = ~({in6[4]} | csa_tree_add_48_2_groupi_n_175);
 assign csa_tree_add_48_2_groupi_n_366 = ~(csa_tree_add_48_2_groupi_n_170 & {in6[3]});
 assign csa_tree_add_48_2_groupi_n_365 = ~({in4[4]} | csa_tree_add_48_2_groupi_n_140);
 assign csa_tree_add_48_2_groupi_n_364 = ~({in4[5]} | csa_tree_add_48_2_groupi_n_167);
 assign csa_tree_add_48_2_groupi_n_363 = ~(csa_tree_add_48_2_groupi_n_137 & {in2[2]});
 assign csa_tree_add_48_2_groupi_n_362 = ~({in2[6]} | csa_tree_add_48_2_groupi_n_136);
 assign csa_tree_add_48_2_groupi_n_361 = ~(csa_tree_add_48_2_groupi_n_168 & {in4[7]});
 assign csa_tree_add_48_2_groupi_n_360 = ~({in4[5]} | csa_tree_add_48_2_groupi_n_168);
 assign csa_tree_add_48_2_groupi_n_359 = ~({in6[4]} | csa_tree_add_48_2_groupi_n_141);
 assign csa_tree_add_48_2_groupi_n_358 = ~({in6[6]} | csa_tree_add_48_2_groupi_n_139);
 assign csa_tree_add_48_2_groupi_n_357 = ~(csa_tree_add_48_2_groupi_n_166 & {in2[5]});
 assign csa_tree_add_48_2_groupi_n_356 = ~(csa_tree_add_48_2_groupi_n_201 & {in6[3]});
 assign csa_tree_add_48_2_groupi_n_355 = ~({in4[2]} | csa_tree_add_48_2_groupi_n_140);
 assign csa_tree_add_48_2_groupi_n_354 = ~({in2[7]} | csa_tree_add_48_2_groupi_n_166);
 assign csa_tree_add_48_2_groupi_n_353 = ~({in4[4]} | csa_tree_add_48_2_groupi_n_174);
 assign csa_tree_add_48_2_groupi_n_352 = ~({in4[3]} | csa_tree_add_48_2_groupi_n_167);
 assign csa_tree_add_48_2_groupi_n_351 = ~({in2[3]} | csa_tree_add_48_2_groupi_n_198);
 assign csa_tree_add_48_2_groupi_n_350 = ~({in4[3]} | csa_tree_add_48_2_groupi_n_199);
 assign csa_tree_add_48_2_groupi_n_349 = ~(csa_tree_add_48_2_groupi_n_173 & {in4[6]});
 assign csa_tree_add_48_2_groupi_n_348 = ~({in2[2]} | csa_tree_add_48_2_groupi_n_171);
 assign csa_tree_add_48_2_groupi_n_347 = ~(csa_tree_add_48_2_groupi_n_175 & {in6[4]});
 assign csa_tree_add_48_2_groupi_n_346 = ~({in6[3]} | csa_tree_add_48_2_groupi_n_170);
 assign csa_tree_add_48_2_groupi_n_345 = ~(csa_tree_add_48_2_groupi_n_196 & {in2[1]});
 assign csa_tree_add_48_2_groupi_n_344 = ~(csa_tree_add_48_2_groupi_n_174 & {in3[4]});
 assign csa_tree_add_48_2_groupi_n_343 = ~(csa_tree_add_48_2_groupi_n_175 & {in5[6]});
 assign csa_tree_add_48_2_groupi_n_342 = ~(csa_tree_add_48_2_groupi_n_177 & {in5[6]});
 assign csa_tree_add_48_2_groupi_n_341 = ~(csa_tree_add_48_2_groupi_n_162 & {in4[3]});
 assign csa_tree_add_48_2_groupi_n_340 = ~(csa_tree_add_48_2_groupi_n_141 & {in5[2]});
 assign csa_tree_add_48_2_groupi_n_339 = ~(csa_tree_add_48_2_groupi_n_173 & {in3[2]});
 assign csa_tree_add_48_2_groupi_n_338 = ~(csa_tree_add_48_2_groupi_n_184 & {in4[5]});
 assign csa_tree_add_48_2_groupi_n_337 = ~(csa_tree_add_48_2_groupi_n_141 & {in5[4]});
 assign csa_tree_add_48_2_groupi_n_336 = ~(csa_tree_add_48_2_groupi_n_140 & {in3[1]});
 assign csa_tree_add_48_2_groupi_n_335 = ~(csa_tree_add_48_2_groupi_n_151 & {in4[5]});
 assign csa_tree_add_48_2_groupi_n_334 = ~(csa_tree_add_48_2_groupi_n_155 & {in6[3]});
 assign csa_tree_add_48_2_groupi_n_415 = ~(csa_tree_add_48_2_groupi_n_163 & {in2[1]});
 assign csa_tree_add_48_2_groupi_n_333 = ~(csa_tree_add_48_2_groupi_n_155 & {in6[5]});
 assign csa_tree_add_48_2_groupi_n_332 = ~({in5[1]} | csa_tree_add_48_2_groupi_n_139);
 assign csa_tree_add_48_2_groupi_n_331 = ~(csa_tree_add_48_2_groupi_n_141 & {in5[5]});
 assign csa_tree_add_48_2_groupi_n_330 = ~({in2[7]} & {in1[23]});
 assign csa_tree_add_48_2_groupi_n_414 = ~({in6[7]} & {in5[1]});
 assign csa_tree_add_48_2_groupi_n_413 = ~({in2[7]} & {in1[1]});
 assign csa_tree_add_48_2_groupi_n_412 = ~({in6[0]} & {in6[1]});
 assign csa_tree_add_48_2_groupi_n_411 = ~({in4[0]} & {in4[1]});
 assign csa_tree_add_48_2_groupi_n_329 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_143);
 assign csa_tree_add_48_2_groupi_n_328 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_148);
 assign csa_tree_add_48_2_groupi_n_327 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_185);
 assign csa_tree_add_48_2_groupi_n_326 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_186);
 assign csa_tree_add_48_2_groupi_n_325 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_163);
 assign csa_tree_add_48_2_groupi_n_324 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_154);
 assign csa_tree_add_48_2_groupi_n_323 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_159);
 assign csa_tree_add_48_2_groupi_n_322 = ~(csa_tree_add_48_2_groupi_n_139 | csa_tree_add_48_2_groupi_n_155);
 assign csa_tree_add_48_2_groupi_n_321 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_150);
 assign csa_tree_add_48_2_groupi_n_320 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_152);
 assign csa_tree_add_48_2_groupi_n_319 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_193);
 assign csa_tree_add_48_2_groupi_n_318 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_164);
 assign csa_tree_add_48_2_groupi_n_317 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_160);
 assign csa_tree_add_48_2_groupi_n_316 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_149);
 assign csa_tree_add_48_2_groupi_n_315 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_157);
 assign csa_tree_add_48_2_groupi_n_314 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_196);
 assign csa_tree_add_48_2_groupi_n_313 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_189);
 assign csa_tree_add_48_2_groupi_n_312 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_195);
 assign csa_tree_add_48_2_groupi_n_410 = ~({in2[7]} & {in1[2]});
 assign csa_tree_add_48_2_groupi_n_311 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_145);
 assign csa_tree_add_48_2_groupi_n_409 = ~({in6[7]} & {in5[2]});
 assign csa_tree_add_48_2_groupi_n_407 = ~({in4[0]} & {in3[0]});
 assign csa_tree_add_48_2_groupi_n_310 = ~(csa_tree_add_48_2_groupi_n_136 | csa_tree_add_48_2_groupi_n_156);
 assign csa_tree_add_48_2_groupi_n_406 = ~({in4[7]} & {in3[3]});
 assign csa_tree_add_48_2_groupi_n_405 = ~({in4[7]} & {in3[2]});
 assign csa_tree_add_48_2_groupi_n_309 = ~(csa_tree_add_48_2_groupi_n_173 | csa_tree_add_48_2_groupi_n_162);
 assign csa_tree_add_48_2_groupi_n_308 = ~(csa_tree_add_48_2_groupi_n_139 | csa_tree_add_48_2_groupi_n_192);
 assign csa_tree_add_48_2_groupi_n_403 = ~({in6[0]} & {in5[0]});
 assign csa_tree_add_48_2_groupi_n_402 = ~({in2[7]} & {in1[7]});
 assign csa_tree_add_48_2_groupi_n_303 = ~(csa_tree_add_48_2_groupi_n_185 & {in2[1]});
 assign csa_tree_add_48_2_groupi_n_302 = ~({in5[5]} | csa_tree_add_48_2_groupi_n_175);
 assign csa_tree_add_48_2_groupi_n_301 = ~(csa_tree_add_48_2_groupi_n_149 & {in2[1]});
 assign csa_tree_add_48_2_groupi_n_300 = ~({in2[1]} | csa_tree_add_48_2_groupi_n_157);
 assign csa_tree_add_48_2_groupi_n_299 = ~(csa_tree_add_48_2_groupi_n_137 & {in1[10]});
 assign csa_tree_add_48_2_groupi_n_298 = ~(csa_tree_add_48_2_groupi_n_194 & {in2[5]});
 assign csa_tree_add_48_2_groupi_n_297 = ~(csa_tree_add_48_2_groupi_n_141 & {in5[7]});
 assign csa_tree_add_48_2_groupi_n_296 = ~(csa_tree_add_48_2_groupi_n_177 & {in5[4]});
 assign csa_tree_add_48_2_groupi_n_295 = ~({in6[1]} | csa_tree_add_48_2_groupi_n_146);
 assign csa_tree_add_48_2_groupi_n_294 = ~({in4[1]} | csa_tree_add_48_2_groupi_n_161);
 assign csa_tree_add_48_2_groupi_n_293 = ~(csa_tree_add_48_2_groupi_n_158 & {in2[1]});
 assign csa_tree_add_48_2_groupi_n_307 = ~(csa_tree_add_48_2_groupi_n_137 & {in1[3]});
 assign csa_tree_add_48_2_groupi_n_292 = ~(csa_tree_add_48_2_groupi_n_158 & {in2[3]});
 assign csa_tree_add_48_2_groupi_n_291 = ~(csa_tree_add_48_2_groupi_n_177 & {in5[7]});
 assign csa_tree_add_48_2_groupi_n_290 = ~(csa_tree_add_48_2_groupi_n_161 & {in4[3]});
 assign csa_tree_add_48_2_groupi_n_289 = ~(csa_tree_add_48_2_groupi_n_158 & {in2[7]});
 assign csa_tree_add_48_2_groupi_n_288 = ~(csa_tree_add_48_2_groupi_n_184 & {in4[1]});
 assign csa_tree_add_48_2_groupi_n_287 = ~({in5[1]} | csa_tree_add_48_2_groupi_n_177);
 assign csa_tree_add_48_2_groupi_n_286 = ~(csa_tree_add_48_2_groupi_n_140 & {in3[6]});
 assign csa_tree_add_48_2_groupi_n_285 = ~(csa_tree_add_48_2_groupi_n_173 & {in3[3]});
 assign csa_tree_add_48_2_groupi_n_284 = ~(csa_tree_add_48_2_groupi_n_187 & {in4[3]});
 assign csa_tree_add_48_2_groupi_n_283 = ~({in5[5]} | csa_tree_add_48_2_groupi_n_177);
 assign csa_tree_add_48_2_groupi_n_282 = ~(csa_tree_add_48_2_groupi_n_192 & {in6[1]});
 assign csa_tree_add_48_2_groupi_n_281 = ~(csa_tree_add_48_2_groupi_n_148 & {in2[1]});
 assign csa_tree_add_48_2_groupi_n_280 = ~(csa_tree_add_48_2_groupi_n_183 & {in6[1]});
 assign csa_tree_add_48_2_groupi_n_279 = ~(csa_tree_add_48_2_groupi_n_174 & {in3[1]});
 assign csa_tree_add_48_2_groupi_n_278 = ~(csa_tree_add_48_2_groupi_n_141 & {in5[6]});
 assign csa_tree_add_48_2_groupi_n_277 = ~({in5[2]} | csa_tree_add_48_2_groupi_n_177);
 assign csa_tree_add_48_2_groupi_n_276 = ~(csa_tree_add_48_2_groupi_n_137 & {in1[11]});
 assign csa_tree_add_48_2_groupi_n_275 = ~({in6[1]} | csa_tree_add_48_2_groupi_n_188);
 assign csa_tree_add_48_2_groupi_n_274 = ~(csa_tree_add_48_2_groupi_n_176 & {in3[2]});
 assign csa_tree_add_48_2_groupi_n_273 = ~(csa_tree_add_48_2_groupi_n_194 & {in2[7]});
 assign csa_tree_add_48_2_groupi_n_272 = ~(csa_tree_add_48_2_groupi_n_190 & {in4[5]});
 assign csa_tree_add_48_2_groupi_n_271 = ~(csa_tree_add_48_2_groupi_n_164 & {in2[1]});
 assign csa_tree_add_48_2_groupi_n_270 = ~({in3[5]} | csa_tree_add_48_2_groupi_n_176);
 assign csa_tree_add_48_2_groupi_n_306 = ~(csa_tree_add_48_2_groupi_n_191 & {in4[1]});
 assign csa_tree_add_48_2_groupi_n_305 = ~(csa_tree_add_48_2_groupi_n_176 & {in3[3]});
 assign csa_tree_add_48_2_groupi_n_269 = ~(csa_tree_add_48_2_groupi_n_188 & {in6[5]});
 assign csa_tree_add_48_2_groupi_n_268 = ~(csa_tree_add_48_2_groupi_n_182 & {in2[3]});
 assign csa_tree_add_48_2_groupi_n_267 = ~(csa_tree_add_48_2_groupi_n_147 & {in6[5]});
 assign csa_tree_add_48_2_groupi_n_266 = ~(csa_tree_add_48_2_groupi_n_136 & {in1[1]});
 assign csa_tree_add_48_2_groupi_n_265 = ~({in1[4]} | csa_tree_add_48_2_groupi_n_137);
 assign csa_tree_add_48_2_groupi_n_264 = ~(csa_tree_add_48_2_groupi_n_147 & {in6[1]});
 assign csa_tree_add_48_2_groupi_n_263 = ~(csa_tree_add_48_2_groupi_n_136 & {in1[2]});
 assign csa_tree_add_48_2_groupi_n_262 = ~(csa_tree_add_48_2_groupi_n_162 & {in4[5]});
 assign csa_tree_add_48_2_groupi_n_261 = ~(csa_tree_add_48_2_groupi_n_174 & {in3[6]});
 assign csa_tree_add_48_2_groupi_n_260 = ~(csa_tree_add_48_2_groupi_n_141 & {in5[1]});
 assign csa_tree_add_48_2_groupi_n_259 = ~({in3[4]} | csa_tree_add_48_2_groupi_n_176);
 assign csa_tree_add_48_2_groupi_n_258 = ~(csa_tree_add_48_2_groupi_n_137 & {in1[5]});
 assign csa_tree_add_48_2_groupi_n_257 = ~(csa_tree_add_48_2_groupi_n_183 & {in6[3]});
 assign csa_tree_add_48_2_groupi_n_256 = ~({in6[3]} | csa_tree_add_48_2_groupi_n_188);
 assign csa_tree_add_48_2_groupi_n_255 = ~(csa_tree_add_48_2_groupi_n_137 & {in1[9]});
 assign csa_tree_add_48_2_groupi_n_254 = ~(csa_tree_add_48_2_groupi_n_140 & {in3[4]});
 assign csa_tree_add_48_2_groupi_n_253 = ~({in5[1]} | csa_tree_add_48_2_groupi_n_175);
 assign csa_tree_add_48_2_groupi_n_252 = ~({in6[7]} | csa_tree_add_48_2_groupi_n_146);
 assign csa_tree_add_48_2_groupi_n_251 = ~(csa_tree_add_48_2_groupi_n_144 & {in6[7]});
 assign csa_tree_add_48_2_groupi_n_250 = ~(csa_tree_add_48_2_groupi_n_161 & {in4[5]});
 assign csa_tree_add_48_2_groupi_n_249 = ~({in4[1]} | csa_tree_add_48_2_groupi_n_190);
 assign csa_tree_add_48_2_groupi_n_248 = ~({in6[3]} | csa_tree_add_48_2_groupi_n_146);
 assign csa_tree_add_48_2_groupi_n_247 = ~(csa_tree_add_48_2_groupi_n_146 & {in6[5]});
 assign csa_tree_add_48_2_groupi_n_246 = ~(csa_tree_add_48_2_groupi_n_138 & {in1[5]});
 assign csa_tree_add_48_2_groupi_n_245 = ~(csa_tree_add_48_2_groupi_n_191 & {in4[7]});
 assign csa_tree_add_48_2_groupi_n_244 = ~(csa_tree_add_48_2_groupi_n_174 & {in3[7]});
 assign csa_tree_add_48_2_groupi_n_243 = ~(csa_tree_add_48_2_groupi_n_148 & {in2[3]});
 assign csa_tree_add_48_2_groupi_n_242 = ~(csa_tree_add_48_2_groupi_n_163 & {in2[7]});
 assign csa_tree_add_48_2_groupi_n_241 = ~(csa_tree_add_48_2_groupi_n_183 & {in6[5]});
 assign csa_tree_add_48_2_groupi_n_240 = ~(csa_tree_add_48_2_groupi_n_174 & {in3[3]});
 assign csa_tree_add_48_2_groupi_n_239 = ~(csa_tree_add_48_2_groupi_n_138 & {in1[1]});
 assign csa_tree_add_48_2_groupi_n_238 = ~(csa_tree_add_48_2_groupi_n_191 & {in4[5]});
 assign csa_tree_add_48_2_groupi_n_237 = ~(csa_tree_add_48_2_groupi_n_141 & {in5[3]});
 assign csa_tree_add_48_2_groupi_n_236 = ~({in4[1]} | csa_tree_add_48_2_groupi_n_151);
 assign csa_tree_add_48_2_groupi_n_235 = ~(csa_tree_add_48_2_groupi_n_184 & {in4[7]});
 assign csa_tree_add_48_2_groupi_n_234 = ~(csa_tree_add_48_2_groupi_n_140 & {in3[5]});
 assign csa_tree_add_48_2_groupi_n_233 = ~(csa_tree_add_48_2_groupi_n_174 & {in3[2]});
 assign csa_tree_add_48_2_groupi_n_232 = ~(csa_tree_add_48_2_groupi_n_192 & {in6[5]});
 assign csa_tree_add_48_2_groupi_n_231 = ~(csa_tree_add_48_2_groupi_n_171 & {in1[2]});
 assign csa_tree_add_48_2_groupi_n_230 = ~(csa_tree_add_48_2_groupi_n_190 & {in4[3]});
 assign csa_tree_add_48_2_groupi_n_229 = ~(csa_tree_add_48_2_groupi_n_187 & {in4[5]});
 assign csa_tree_add_48_2_groupi_n_228 = ~(csa_tree_add_48_2_groupi_n_177 & {in5[3]});
 assign csa_tree_add_48_2_groupi_n_227 = ~(csa_tree_add_48_2_groupi_n_144 & {in6[5]});
 assign csa_tree_add_48_2_groupi_n_226 = ~({in3[1]} | csa_tree_add_48_2_groupi_n_176);
 assign csa_tree_add_48_2_groupi_n_225 = ~(csa_tree_add_48_2_groupi_n_175 & {in5[4]});
 assign csa_tree_add_48_2_groupi_n_224 = ~(csa_tree_add_48_2_groupi_n_137 & {in1[2]});
 assign csa_tree_add_48_2_groupi_n_223 = ~(csa_tree_add_48_2_groupi_n_171 & {in1[7]});
 assign csa_tree_add_48_2_groupi_n_222 = ~(csa_tree_add_48_2_groupi_n_149 & {in2[5]});
 assign csa_tree_add_48_2_groupi_n_221 = ~(csa_tree_add_48_2_groupi_n_137 & {in1[1]});
 assign csa_tree_add_48_2_groupi_n_220 = ~(csa_tree_add_48_2_groupi_n_151 & {in4[3]});
 assign csa_tree_add_48_2_groupi_n_219 = ~({in3[6]} | csa_tree_add_48_2_groupi_n_176);
 assign csa_tree_add_48_2_groupi_n_216 = ~({in5[0]} | csa_tree_add_48_2_groupi_n_139);
 assign csa_tree_add_48_2_groupi_n_211 = ~(csa_tree_add_48_2_groupi_n_180 & {in6[3]});
 assign csa_tree_add_48_2_groupi_n_210 = ~({in6[7]} | csa_tree_add_48_2_groupi_n_180);
 assign csa_tree_add_48_2_groupi_n_209 = ~(csa_tree_add_48_2_groupi_n_178 & {in4[3]});
 assign csa_tree_add_48_2_groupi_n_208 = ~(csa_tree_add_48_2_groupi_n_140 & {in3[0]});
 assign csa_tree_add_48_2_groupi_n_207 = ~(csa_tree_add_48_2_groupi_n_175 & {in5[0]});
 assign csa_tree_add_48_2_groupi_n_206 = ~(csa_tree_add_48_2_groupi_n_141 & {in5[0]});
 assign csa_tree_add_48_2_groupi_n_205 = ~(csa_tree_add_48_2_groupi_n_180 & {in6[5]});
 assign csa_tree_add_48_2_groupi_n_204 = ~(csa_tree_add_48_2_groupi_n_179 & {in2[7]});
 assign csa_tree_add_48_2_groupi_n_203 = ~(csa_tree_add_48_2_groupi_n_136 & {in1[0]});
 assign csa_tree_add_48_2_groupi_n_304 = ~({in2[0]} & {in2[1]});
 assign csa_tree_add_48_2_groupi_n_202 = ({in4[7]} & {in3[0]});
 assign csa_tree_add_48_2_groupi_n_201 = ~{in6[2]};
 assign csa_tree_add_48_2_groupi_n_200 = ~{in6[6]};
 assign csa_tree_add_48_2_groupi_n_199 = ~{in4[2]};
 assign csa_tree_add_48_2_groupi_n_198 = ~{in2[2]};
 assign csa_tree_add_48_2_groupi_n_197 = ~{in1[25]};
 assign csa_tree_add_48_2_groupi_n_196 = ~{in1[11]};
 assign csa_tree_add_48_2_groupi_n_195 = ~{in1[13]};
 assign csa_tree_add_48_2_groupi_n_194 = ~{in1[1]};
 assign csa_tree_add_48_2_groupi_n_193 = ~{in1[20]};
 assign csa_tree_add_48_2_groupi_n_192 = ~{in5[3]};
 assign csa_tree_add_48_2_groupi_n_191 = ~{in3[3]};
 assign csa_tree_add_48_2_groupi_n_190 = ~{in3[6]};
 assign csa_tree_add_48_2_groupi_n_189 = ~{in1[6]};
 assign csa_tree_add_48_2_groupi_n_188 = ~{in5[5]};
 assign csa_tree_add_48_2_groupi_n_187 = ~{in3[7]};
 assign csa_tree_add_48_2_groupi_n_186 = ~{in1[12]};
 assign csa_tree_add_48_2_groupi_n_185 = ~{in1[10]};
 assign csa_tree_add_48_2_groupi_n_184 = ~{in3[2]};
 assign csa_tree_add_48_2_groupi_n_183 = ~{in5[7]};
 assign csa_tree_add_48_2_groupi_n_182 = ~{in1[7]};
 assign csa_tree_add_48_2_groupi_n_181 = ~{in4[0]};
 assign csa_tree_add_48_2_groupi_n_180 = ~{in5[0]};
 assign csa_tree_add_48_2_groupi_n_179 = ~{in1[0]};
 assign csa_tree_add_48_2_groupi_n_178 = ~{in3[0]};
 assign csa_tree_add_48_2_groupi_n_177 = ~{in6[1]};
 assign csa_tree_add_48_2_groupi_n_176 = ~{in4[1]};
 assign csa_tree_add_48_2_groupi_n_175 = ~{in6[3]};
 assign csa_tree_add_48_2_groupi_n_174 = ~{in4[5]};
 assign csa_tree_add_48_2_groupi_n_173 = ~{in4[7]};
 assign csa_tree_add_48_2_groupi_n_172 = ~{in2[0]};
 assign csa_tree_add_48_2_groupi_n_171 = ~{in2[3]};
 assign csa_tree_add_48_2_groupi_n_170 = ~{in6[4]};
 assign csa_tree_add_48_2_groupi_n_169 = ~{in2[4]};
 assign csa_tree_add_48_2_groupi_n_168 = ~{in4[6]};
 assign csa_tree_add_48_2_groupi_n_167 = ~{in4[4]};
 assign csa_tree_add_48_2_groupi_n_166 = ~{in2[6]};
 assign csa_tree_add_48_2_groupi_n_165 = ~{in1[24]};
 assign csa_tree_add_48_2_groupi_n_164 = ~{in1[14]};
 assign csa_tree_add_48_2_groupi_n_163 = ~{in1[3]};
 assign csa_tree_add_48_2_groupi_n_162 = ~{in3[1]};
 assign csa_tree_add_48_2_groupi_n_161 = ~{in3[5]};
 assign csa_tree_add_48_2_groupi_n_160 = ~{in1[21]};
 assign csa_tree_add_48_2_groupi_n_159 = ~{in1[19]};
 assign csa_tree_add_48_2_groupi_n_158 = ~{in1[2]};
 assign csa_tree_add_48_2_groupi_n_157 = ~{in1[4]};
 assign csa_tree_add_48_2_groupi_n_156 = ~{in1[15]};
 assign csa_tree_add_48_2_groupi_n_155 = ~{in5[4]};
 assign csa_tree_add_48_2_groupi_n_154 = ~{in1[17]};
 assign csa_tree_add_48_2_groupi_n_153 = ~{in1[23]};
 assign csa_tree_add_48_2_groupi_n_152 = ~{in1[16]};
 assign csa_tree_add_48_2_groupi_n_151 = ~{in3[4]};
 assign csa_tree_add_48_2_groupi_n_150 = ~{in1[18]};
 assign csa_tree_add_48_2_groupi_n_149 = ~{in1[5]};
 assign csa_tree_add_48_2_groupi_n_148 = ~{in1[9]};
 assign csa_tree_add_48_2_groupi_n_147 = ~{in5[6]};
 assign csa_tree_add_48_2_groupi_n_146 = ~{in5[1]};
 assign csa_tree_add_48_2_groupi_n_145 = ~{in1[22]};
 assign csa_tree_add_48_2_groupi_n_144 = ~{in5[2]};
 assign csa_tree_add_48_2_groupi_n_143 = ~{in1[8]};
 assign csa_tree_add_48_2_groupi_n_142 = ~{in6[0]};
 assign csa_tree_add_48_2_groupi_n_141 = ~{in6[5]};
 assign csa_tree_add_48_2_groupi_n_140 = ~{in4[3]};
 assign csa_tree_add_48_2_groupi_n_139 = ~{in6[7]};
 assign csa_tree_add_48_2_groupi_n_138 = ~{in2[5]};
 assign csa_tree_add_48_2_groupi_n_137 = ~{in2[1]};
 assign csa_tree_add_48_2_groupi_n_136 = ~{in2[7]};
 assign csa_tree_add_48_2_groupi_n_114 = ({in6[7]} & {in5[0]});
 assign csa_tree_add_48_2_groupi_n_113 = ({in6[6]} | {in5[0]});
 assign csa_tree_add_48_2_groupi_n_112 = ({in2[6]} | {in1[0]});
 assign csa_tree_add_48_2_groupi_n_111 = ({in2[4]} | {in1[0]});
 assign csa_tree_add_48_2_groupi_n_110 = ({in4[6]} | {in3[0]});
 assign csa_tree_add_48_2_groupi_n_109 = ({in2[0]} & {in1[0]});
 assign csa_tree_add_48_2_groupi_n_107 = (csa_tree_add_48_2_groupi_n_1718 ^ csa_tree_add_48_2_groupi_n_1673);
 assign csa_tree_add_48_2_groupi_n_106 = (csa_tree_add_48_2_groupi_n_1678 & csa_tree_add_48_2_groupi_n_1665);
 assign csa_tree_add_48_2_groupi_n_104 = ~(csa_tree_add_48_2_groupi_n_1650 ^ n_164);
 assign csa_tree_add_48_2_groupi_n_103 = (csa_tree_add_48_2_groupi_n_101 ^ csa_tree_add_48_2_groupi_n_1653);
 assign csa_tree_add_48_2_groupi_n_101 = (csa_tree_add_48_2_groupi_n_1649 ^ csa_tree_add_48_2_groupi_n_1635);
 assign csa_tree_add_48_2_groupi_n_100 = (csa_tree_add_48_2_groupi_n_1594 & csa_tree_add_48_2_groupi_n_1516);
 assign csa_tree_add_48_2_groupi_n_99 = (n_165 ^ csa_tree_add_48_2_groupi_n_1591);
 assign csa_tree_add_48_2_groupi_n_97 = (csa_tree_add_48_2_groupi_n_87 | csa_tree_add_48_2_groupi_n_1536);
 assign csa_tree_add_48_2_groupi_n_96 = (n_169 & csa_tree_add_48_2_groupi_n_1469);
 assign csa_tree_add_48_2_groupi_n_95 = ~(csa_tree_add_48_2_groupi_n_1517 ^ csa_tree_add_48_2_groupi_n_1498);
 assign csa_tree_add_48_2_groupi_n_93 = (csa_tree_add_48_2_groupi_n_85 ^ csa_tree_add_48_2_groupi_n_1519);
 assign csa_tree_add_48_2_groupi_n_92 = ~(csa_tree_add_48_2_groupi_n_1494 ^ csa_tree_add_48_2_groupi_n_1508);
 assign csa_tree_add_48_2_groupi_n_91 = (csa_tree_add_48_2_groupi_n_88 ^ csa_tree_add_48_2_groupi_n_1414);
 assign csa_tree_add_48_2_groupi_n_90 = (csa_tree_add_48_2_groupi_n_1470 & csa_tree_add_48_2_groupi_n_75);
 assign csa_tree_add_48_2_groupi_n_89 = (csa_tree_add_48_2_groupi_n_79 ^ n_171);
 assign csa_tree_add_48_2_groupi_n_88 = (n_172 ^ csa_tree_add_48_2_groupi_n_1417);
 assign csa_tree_add_48_2_groupi_n_87 = (csa_tree_add_48_2_groupi_n_1453 ^ csa_tree_add_48_2_groupi_n_1366);
 assign csa_tree_add_48_2_groupi_n_86 = (csa_tree_add_48_2_groupi_n_72 | csa_tree_add_48_2_groupi_n_1378);
 assign csa_tree_add_48_2_groupi_n_85 = (csa_tree_add_48_2_groupi_n_1474 ^ csa_tree_add_48_2_groupi_n_1408);
 assign csa_tree_add_48_2_groupi_n_84 = (csa_tree_add_48_2_groupi_n_1501 ^ csa_tree_add_48_2_groupi_n_1406);
 assign csa_tree_add_48_2_groupi_n_83 = ~(csa_tree_add_48_2_groupi_n_1377 & ~n_175);
 assign csa_tree_add_48_2_groupi_n_82 = ~(csa_tree_add_48_2_groupi_n_1392 | ~csa_tree_add_48_2_groupi_n_1345);
 assign csa_tree_add_48_2_groupi_n_81 = (n_174 ^ csa_tree_add_48_2_groupi_n_1311);
 assign csa_tree_add_48_2_groupi_n_79 = (csa_tree_add_48_2_groupi_n_1374 ^ csa_tree_add_48_2_groupi_n_1316);
 assign csa_tree_add_48_2_groupi_n_78 = (csa_tree_add_48_2_groupi_n_37 | csa_tree_add_48_2_groupi_n_1191);
 assign csa_tree_add_48_2_groupi_n_77 = ~(csa_tree_add_48_2_groupi_n_1276 ^ csa_tree_add_48_2_groupi_n_1313);
 assign csa_tree_add_48_2_groupi_n_76 = ~(n_174 & ~csa_tree_add_48_2_groupi_n_1311);
 assign csa_tree_add_48_2_groupi_n_75 = ~(csa_tree_add_48_2_groupi_n_55 ^ csa_tree_add_48_2_groupi_n_1310);
 assign csa_tree_add_48_2_groupi_n_74 = ~(csa_tree_add_48_2_groupi_n_1152 ^ csa_tree_add_48_2_groupi_n_1268);
 assign csa_tree_add_48_2_groupi_n_73 = ~(csa_tree_add_48_2_groupi_n_38 & ~csa_tree_add_48_2_groupi_n_1308);
 assign csa_tree_add_48_2_groupi_n_72 = ~(csa_tree_add_48_2_groupi_n_62 ^ csa_tree_add_48_2_groupi_n_1193);
 assign csa_tree_add_48_2_groupi_n_71 = ~(csa_tree_add_48_2_groupi_n_1308 & ~csa_tree_add_48_2_groupi_n_38);
 assign csa_tree_add_48_2_groupi_n_70 = (csa_tree_add_48_2_groupi_n_1284 ^ csa_tree_add_48_2_groupi_n_1197);
 assign csa_tree_add_48_2_groupi_n_65 = (csa_tree_add_48_2_groupi_n_1349 ^ csa_tree_add_48_2_groupi_n_35);
 assign csa_tree_add_48_2_groupi_n_64 = (csa_tree_add_48_2_groupi_n_1273 | csa_tree_add_48_2_groupi_n_1274);
 assign csa_tree_add_48_2_groupi_n_62 = ~(csa_tree_add_48_2_groupi_n_23 ^ csa_tree_add_48_2_groupi_n_1135);
 assign csa_tree_add_48_2_groupi_n_61 = (csa_tree_add_48_2_groupi_n_134 | csa_tree_add_48_2_groupi_n_1360);
 assign csa_tree_add_48_2_groupi_n_60 = ~(csa_tree_add_48_2_groupi_n_132 | ~csa_tree_add_48_2_groupi_n_1115);
 assign csa_tree_add_48_2_groupi_n_55 = ~(n_180 ^ csa_tree_add_48_2_groupi_n_1124);
 assign csa_tree_add_48_2_groupi_n_53 = (csa_tree_add_48_2_groupi_n_51 ^ csa_tree_add_48_2_groupi_n_1086);
 assign csa_tree_add_48_2_groupi_n_52 = ~(csa_tree_add_48_2_groupi_n_1082 ^ csa_tree_add_48_2_groupi_n_1083);
 assign csa_tree_add_48_2_groupi_n_51 = ~(csa_tree_add_48_2_groupi_n_1005 ^ csa_tree_add_48_2_groupi_n_1073);
 assign csa_tree_add_48_2_groupi_n_50 = ~(csa_tree_add_48_2_groupi_n_52 ^ csa_tree_add_48_2_groupi_n_1050);
 assign csa_tree_add_48_2_groupi_n_49 = ~(csa_tree_add_48_2_groupi_n_1078 | ~csa_tree_add_48_2_groupi_n_130);
 assign csa_tree_add_48_2_groupi_n_46 = ~(csa_tree_add_48_2_groupi_n_1118 ^ csa_tree_add_48_2_groupi_n_1015);
 assign csa_tree_add_48_2_groupi_n_45 = (csa_tree_add_48_2_groupi_n_1008 ^ csa_tree_add_48_2_groupi_n_1010);
 assign csa_tree_add_48_2_groupi_n_44 = ~(csa_tree_add_48_2_groupi_n_1074 | ~csa_tree_add_48_2_groupi_n_1007);
 assign csa_tree_add_48_2_groupi_n_43 = ~(csa_tree_add_48_2_groupi_n_1071 | ~csa_tree_add_48_2_groupi_n_1006);
 assign csa_tree_add_48_2_groupi_n_41 = ~(csa_tree_add_48_2_groupi_n_28 | ~csa_tree_add_48_2_groupi_n_1003);
 assign csa_tree_add_48_2_groupi_n_40 = ~(csa_tree_add_48_2_groupi_n_1080 | ~csa_tree_add_48_2_groupi_n_1002);
 assign csa_tree_add_48_2_groupi_n_39 = ~(csa_tree_add_48_2_groupi_n_405 | ~csa_tree_add_48_2_groupi_n_1000);
 assign csa_tree_add_48_2_groupi_n_38 = (csa_tree_add_48_2_groupi_n_1119 ^ csa_tree_add_48_2_groupi_n_944);
 assign csa_tree_add_48_2_groupi_n_37 = ~(csa_tree_add_48_2_groupi_n_1092 ^ csa_tree_add_48_2_groupi_n_943);
 assign csa_tree_add_48_2_groupi_n_35 = ~(csa_tree_add_48_2_groupi_n_45 ^ csa_tree_add_48_2_groupi_n_937);
 assign csa_tree_add_48_2_groupi_n_31 = ~(csa_tree_add_48_2_groupi_n_681 & ~csa_tree_add_48_2_groupi_n_584);
 assign csa_tree_add_48_2_groupi_n_30 = ~(csa_tree_add_48_2_groupi_n_553 | ~csa_tree_add_48_2_groupi_n_751);
 assign csa_tree_add_48_2_groupi_n_29 = ~(csa_tree_add_48_2_groupi_n_723 | ~csa_tree_add_48_2_groupi_n_494);
 assign csa_tree_add_48_2_groupi_n_28 = ~(csa_tree_add_48_2_groupi_n_993 | ~csa_tree_add_48_2_groupi_n_748);
 assign csa_tree_add_48_2_groupi_n_27 = ~(csa_tree_add_48_2_groupi_n_844 & ~csa_tree_add_48_2_groupi_n_747);
 assign csa_tree_add_48_2_groupi_n_26 = ~(csa_tree_add_48_2_groupi_n_830 | ~csa_tree_add_48_2_groupi_n_746);
 assign csa_tree_add_48_2_groupi_n_25 = ~(csa_tree_add_48_2_groupi_n_802 & ~csa_tree_add_48_2_groupi_n_745);
 assign csa_tree_add_48_2_groupi_n_24 = (csa_tree_add_48_2_groupi_n_744 & (csa_tree_add_48_2_groupi_n_726
    | csa_tree_add_48_2_groupi_n_140));
 assign csa_tree_add_48_2_groupi_n_23 = ~(csa_tree_add_48_2_groupi_n_982 ^ csa_tree_add_48_2_groupi_n_734);
 assign csa_tree_add_48_2_groupi_n_22 = ~(csa_tree_add_48_2_groupi_n_981 ^ csa_tree_add_48_2_groupi_n_731);
 assign csa_tree_add_48_2_groupi_n_21 = ~(csa_tree_add_48_2_groupi_n_141 | ~csa_tree_add_48_2_groupi_n_728);
 assign csa_tree_add_48_2_groupi_n_20 = ~(csa_tree_add_48_2_groupi_n_444 | ~csa_tree_add_48_2_groupi_n_678);
 assign csa_tree_add_48_2_groupi_n_19 = ~(csa_tree_add_48_2_groupi_n_121 & ~csa_tree_add_48_2_groupi_n_605);
 assign csa_tree_add_48_2_groupi_n_18 = ~(n_189 & ~csa_tree_add_48_2_groupi_n_558);
 assign csa_tree_add_48_2_groupi_n_17 = (csa_tree_add_48_2_groupi_n_555 ^ csa_tree_add_48_2_groupi_n_554);
 assign csa_tree_add_48_2_groupi_n_16 = ~(csa_tree_add_48_2_groupi_n_470 | ~csa_tree_add_48_2_groupi_n_551);
 assign csa_tree_add_48_2_groupi_n_15 = ~(csa_tree_add_48_2_groupi_n_123 & ~csa_tree_add_48_2_groupi_n_518);
 assign csa_tree_add_48_2_groupi_n_14 = ~(csa_tree_add_48_2_groupi_n_543 | ~csa_tree_add_48_2_groupi_n_517);
 assign csa_tree_add_48_2_groupi_n_13 = ~(csa_tree_add_48_2_groupi_n_124 | ~csa_tree_add_48_2_groupi_n_514);
 assign csa_tree_add_48_2_groupi_n_12 = ~(csa_tree_add_48_2_groupi_n_543 | ~csa_tree_add_48_2_groupi_n_511);
 assign csa_tree_add_48_2_groupi_n_11 = ~(csa_tree_add_48_2_groupi_n_544 & ~csa_tree_add_48_2_groupi_n_508);
 assign csa_tree_add_48_2_groupi_n_10 = ~({in6[0]} & ~csa_tree_add_48_2_groupi_n_490);
 assign csa_tree_add_48_2_groupi_n_9 = ~({in4[0]} & ~csa_tree_add_48_2_groupi_n_489);
 assign csa_tree_add_48_2_groupi_n_8 = ~(csa_tree_add_48_2_groupi_n_729 | ~csa_tree_add_48_2_groupi_n_481);
 assign csa_tree_add_48_2_groupi_n_7 = ~(csa_tree_add_48_2_groupi_n_727 & ~csa_tree_add_48_2_groupi_n_470);
 assign csa_tree_add_48_2_groupi_n_6 = ~(csa_tree_add_48_2_groupi_n_126 | ~csa_tree_add_48_2_groupi_n_468);
 assign csa_tree_add_48_2_groupi_n_5 = ~(csa_tree_add_48_2_groupi_n_118 | ~csa_tree_add_48_2_groupi_n_467);
 assign csa_tree_add_48_2_groupi_n_4 = ~(csa_tree_add_48_2_groupi_n_551 & ~csa_tree_add_48_2_groupi_n_466);
 assign csa_tree_add_48_2_groupi_n_3 = ~(csa_tree_add_48_2_groupi_n_722 | ~csa_tree_add_48_2_groupi_n_465);
 assign csa_tree_add_48_2_groupi_n_2 = ~(csa_tree_add_48_2_groupi_n_541 | ~csa_tree_add_48_2_groupi_n_443);
 assign csa_tree_add_48_2_groupi_n_1 = ~(csa_tree_add_48_2_groupi_n_442 | ~csa_tree_add_48_2_groupi_n_121);
 assign csa_tree_add_48_2_groupi_n_0 = ~(csa_tree_add_48_2_groupi_n_122 | ~csa_tree_add_48_2_groupi_n_434);
 assign csa_tree_add_48_2_groupi_n_134 = (csa_tree_add_48_2_groupi_n_1000 ^ (csa_tree_add_48_2_groupi_n_1018
    ^ csa_tree_add_48_2_groupi_n_405));
 assign {out1[31]} = ~(n_12 ^ n_11);
 assign n_12 = ((n_10 & n_13) | ((n_13 & n_8) | (n_8 & n_10)));
 assign {out1[30]} = (n_13 ^ (n_8 ^ n_10));
 assign n_13 = ((n_9 & n_14) | ((n_14 & n_6) | (n_6 & n_9)));
 assign {out1[29]} = (n_14 ^ (n_6 ^ n_9));
 assign n_14 = ((n_7 & n_15) | ((n_15 & n_4) | (n_4 & n_7)));
 assign {out1[28]} = (n_15 ^ (n_4 ^ n_7));
 assign n_15 = ((n_5 & n_16) | ((n_16 & n_2) | (n_2 & n_5)));
 assign {out1[27]} = (n_16 ^ (n_2 ^ n_5));
 assign n_16 = ((n_0 & n_3) | ((n_3 & n_1) | (n_1 & n_0)));
 assign {out1[26]} = (n_3 ^ (n_1 ^ n_0));
 assign n_18 = ((csa_tree_add_48_2_groupi_n_1572 & n_20) | ((n_20 & n_28) | (n_28 & csa_tree_add_48_2_groupi_n_1572)));
 assign n_17 = (n_20 ^ (n_28 ^ csa_tree_add_48_2_groupi_n_1572));
 assign n_20 = ((csa_tree_add_48_2_groupi_n_1573 & n_24) | ((n_24 & csa_tree_add_48_2_groupi_n_1564)
    | (csa_tree_add_48_2_groupi_n_1564 & csa_tree_add_48_2_groupi_n_1573)));
 assign n_19 = (n_24 ^ (csa_tree_add_48_2_groupi_n_1564 ^ csa_tree_add_48_2_groupi_n_1573));
 assign n_21 = ~(csa_tree_add_48_2_groupi_n_81 ^ csa_tree_add_48_2_groupi_n_1452);
 assign csa_tree_add_48_2_groupi_n_1452 = ((csa_tree_add_48_2_groupi_n_1089 & csa_tree_add_48_2_groupi_n_50)
    | ((csa_tree_add_48_2_groupi_n_50 & n_35) | (n_35 & csa_tree_add_48_2_groupi_n_1089)));
 assign n_22 = (csa_tree_add_48_2_groupi_n_50 ^ (n_35 ^ csa_tree_add_48_2_groupi_n_1089));
 assign n_24 = ((csa_tree_add_48_2_groupi_n_1565 & n_41) | ((n_41 & csa_tree_add_48_2_groupi_n_1560)
    | (csa_tree_add_48_2_groupi_n_1560 & csa_tree_add_48_2_groupi_n_1565)));
 assign n_23 = (n_41 ^ (csa_tree_add_48_2_groupi_n_1560 ^ csa_tree_add_48_2_groupi_n_1565));
 assign n_25 = ~(csa_tree_add_48_2_groupi_n_1500 ^ n_31);
 assign n_41 = ((csa_tree_add_48_2_groupi_n_1561 & csa_tree_add_48_2_groupi_n_1779) | ((csa_tree_add_48_2_groupi_n_1779
    & csa_tree_add_48_2_groupi_n_1557) | (csa_tree_add_48_2_groupi_n_1557 & csa_tree_add_48_2_groupi_n_1561)));
 assign n_40 = (csa_tree_add_48_2_groupi_n_1779 ^ (csa_tree_add_48_2_groupi_n_1557 ^ csa_tree_add_48_2_groupi_n_1561));
 assign n_37 = ((csa_tree_add_48_2_groupi_n_1433 & csa_tree_add_48_2_groupi_n_1441) | ((csa_tree_add_48_2_groupi_n_1441
    & csa_tree_add_48_2_groupi_n_1212) | (csa_tree_add_48_2_groupi_n_1212 & csa_tree_add_48_2_groupi_n_1433)));
 assign n_36 = (csa_tree_add_48_2_groupi_n_1441 ^ (csa_tree_add_48_2_groupi_n_1212 ^ csa_tree_add_48_2_groupi_n_1433));
 assign n_39 = ((csa_tree_add_48_2_groupi_n_1448 & csa_tree_add_48_2_groupi_n_1432) | ((csa_tree_add_48_2_groupi_n_1432
    & csa_tree_add_48_2_groupi_n_1262) | (csa_tree_add_48_2_groupi_n_1262 & csa_tree_add_48_2_groupi_n_1448)));
 assign n_38 = (csa_tree_add_48_2_groupi_n_1432 ^ (csa_tree_add_48_2_groupi_n_1262 ^ csa_tree_add_48_2_groupi_n_1448));
 assign n_31 = ((csa_tree_add_48_2_groupi_n_1429 & csa_tree_add_48_2_groupi_n_1463) | ((csa_tree_add_48_2_groupi_n_1463
    & csa_tree_add_48_2_groupi_n_1180) | (csa_tree_add_48_2_groupi_n_1180 & csa_tree_add_48_2_groupi_n_1429)));
 assign n_30 = (csa_tree_add_48_2_groupi_n_1463 ^ (csa_tree_add_48_2_groupi_n_1180 ^ csa_tree_add_48_2_groupi_n_1429));
 assign n_27 = ((csa_tree_add_48_2_groupi_n_1431 & csa_tree_add_48_2_groupi_n_1430) | ((csa_tree_add_48_2_groupi_n_1430
    & csa_tree_add_48_2_groupi_n_1258) | (csa_tree_add_48_2_groupi_n_1258 & csa_tree_add_48_2_groupi_n_1431)));
 assign n_26 = (csa_tree_add_48_2_groupi_n_1430 ^ (csa_tree_add_48_2_groupi_n_1258 ^ csa_tree_add_48_2_groupi_n_1431));
 assign n_35 = ((csa_tree_add_48_2_groupi_n_404 & csa_tree_add_48_2_groupi_n_109) | ((csa_tree_add_48_2_groupi_n_109
    & csa_tree_add_48_2_groupi_n_408) | (csa_tree_add_48_2_groupi_n_408 & csa_tree_add_48_2_groupi_n_404)));
 assign n_34 = (csa_tree_add_48_2_groupi_n_109 ^ (csa_tree_add_48_2_groupi_n_408 ^ csa_tree_add_48_2_groupi_n_404));
 assign n_33 = ((csa_tree_add_48_2_groupi_n_1440 & csa_tree_add_48_2_groupi_n_1449) | ((csa_tree_add_48_2_groupi_n_1449
    & csa_tree_add_48_2_groupi_n_1235) | (csa_tree_add_48_2_groupi_n_1235 & csa_tree_add_48_2_groupi_n_1440)));
 assign n_32 = (csa_tree_add_48_2_groupi_n_1449 ^ (csa_tree_add_48_2_groupi_n_1235 ^ csa_tree_add_48_2_groupi_n_1440));
 assign n_29 = ((csa_tree_add_48_2_groupi_n_1423 & csa_tree_add_48_2_groupi_n_1434) | ((csa_tree_add_48_2_groupi_n_1434
    & csa_tree_add_48_2_groupi_n_1254) | (csa_tree_add_48_2_groupi_n_1254 & csa_tree_add_48_2_groupi_n_1423)));
 assign n_28 = (csa_tree_add_48_2_groupi_n_1434 ^ (csa_tree_add_48_2_groupi_n_1254 ^ csa_tree_add_48_2_groupi_n_1423));
 assign n_53 = ~(csa_tree_add_48_2_groupi_n_1755 ^ csa_tree_add_48_2_groupi_n_1710);
 assign n_47 = ~(csa_tree_add_48_2_groupi_n_1774 ^ csa_tree_add_48_2_groupi_n_1620);
 assign n_54 = ~(csa_tree_add_48_2_groupi_n_1770 ^ csa_tree_add_48_2_groupi_n_1667);
 assign n_49 = ~(csa_tree_add_48_2_groupi_n_1766 ^ csa_tree_add_48_2_groupi_n_1697);
 assign n_48 = ~(csa_tree_add_48_2_groupi_n_1763 ^ csa_tree_add_48_2_groupi_n_1696);
 assign n_43 = ~(csa_tree_add_48_2_groupi_n_1759 ^ csa_tree_add_48_2_groupi_n_1711);
 assign n_44 = ~(csa_tree_add_48_2_groupi_n_1777 ^ csa_tree_add_48_2_groupi_n_1613);
 assign n_45 = ~(csa_tree_add_48_2_groupi_n_1704 ^ csa_tree_add_48_2_groupi_n_1655);
 assign n_46 = ~(csa_tree_add_48_2_groupi_n_1747 ^ csa_tree_add_48_2_groupi_n_1732);
 assign n_42 = ~(csa_tree_add_48_2_groupi_n_1721 ^ csa_tree_add_48_2_groupi_n_1741);
 assign n_55 = ~(csa_tree_add_48_2_groupi_n_1737 ^ csa_tree_add_48_2_groupi_n_1709);
 assign n_50 = ~(csa_tree_add_48_2_groupi_n_1695 ^ csa_tree_add_48_2_groupi_n_1733);
 assign n_51 = ~(csa_tree_add_48_2_groupi_n_1724 ^ csa_tree_add_48_2_groupi_n_1671);
 assign n_52 = ~(csa_tree_add_48_2_groupi_n_1751 ^ csa_tree_add_48_2_groupi_n_1722);
 assign n_57 = ~csa_tree_add_48_2_groupi_n_1625;
 assign n_58 = ~csa_tree_add_48_2_groupi_n_1657;
 assign n_59 = ~csa_tree_add_48_2_groupi_n_1543;
 assign n_56 = ~csa_tree_add_48_2_groupi_n_107;
 assign n_60 = ~csa_tree_add_48_2_groupi_n_1499;
 assign n_164 = (csa_tree_add_48_2_groupi_n_1584 ^ csa_tree_add_48_2_groupi_n_1615);
 assign n_165 = (csa_tree_add_48_2_groupi_n_93 ^ csa_tree_add_48_2_groupi_n_1633);
 assign n_166 = (csa_tree_add_48_2_groupi_n_1614 ^ csa_tree_add_48_2_groupi_n_1601);
 assign n_167 = ~(csa_tree_add_48_2_groupi_n_1592 ^ csa_tree_add_48_2_groupi_n_1523);
 assign n_168 = ~(csa_tree_add_48_2_groupi_n_1544 ^ csa_tree_add_48_2_groupi_n_1537);
 assign n_169 = ~(csa_tree_add_48_2_groupi_n_1490 ^ csa_tree_add_48_2_groupi_n_1387);
 assign n_170 = ~(csa_tree_add_48_2_groupi_n_1450 ^ csa_tree_add_48_2_groupi_n_1345);
 assign n_171 = ~(csa_tree_add_48_2_groupi_n_1340 ^ csa_tree_add_48_2_groupi_n_1280);
 assign n_172 = (csa_tree_add_48_2_groupi_n_1359 ^ csa_tree_add_48_2_groupi_n_1315);
 assign n_173 = (csa_tree_add_48_2_groupi_n_1283 ^ csa_tree_add_48_2_groupi_n_1307);
 assign n_174 = ~(csa_tree_add_48_2_groupi_n_1154 ^ csa_tree_add_48_2_groupi_n_135);
 assign n_175 = (csa_tree_add_48_2_groupi_n_1270 ^ csa_tree_add_48_2_groupi_n_1275);
 assign n_176 = ~(csa_tree_add_48_2_groupi_n_1153 ^ n_177);
 assign n_177 = ~(csa_tree_add_48_2_groupi_n_133 ^ csa_tree_add_48_2_groupi_n_1142);
 assign n_178 = ~(n_181 ^ csa_tree_add_48_2_groupi_n_1016);
 assign n_179 = ~(csa_tree_add_48_2_groupi_n_1116 ^ csa_tree_add_48_2_groupi_n_941);
 assign n_180 = ~(n_183 ^ csa_tree_add_48_2_groupi_n_129);
 assign n_181 = ((csa_tree_add_48_2_groupi_n_1084 & ~csa_tree_add_48_2_groupi_n_1004) | (csa_tree_add_48_2_groupi_n_1085
    & csa_tree_add_48_2_groupi_n_1004));
 assign n_182 = (csa_tree_add_48_2_groupi_n_1019 ^ csa_tree_add_48_2_groupi_n_1020);
 assign n_183 = ~(csa_tree_add_48_2_groupi_n_850 ^ csa_tree_add_48_2_groupi_n_851);
 assign n_185 = ~({in4[0]} | n_184);
 assign n_184 = (csa_tree_add_48_2_groupi_n_176 & ({in4[1]} | csa_tree_add_48_2_groupi_n_181));
 assign n_187 = ~({in6[0]} | n_186);
 assign n_186 = (csa_tree_add_48_2_groupi_n_177 & ({in6[1]} | csa_tree_add_48_2_groupi_n_142));
 assign n_189 = ~({in2[0]} | n_188);
 assign n_188 = (csa_tree_add_48_2_groupi_n_137 & ({in2[1]} | csa_tree_add_48_2_groupi_n_172));
endmodule
