`timescale 1ps / 1ps
module dut_Add2Mul2u8u8u32_4(
          in3,
          in2,
          in1,
          out1,
          clk
);
   input [31:0] in3;
   input [7:0] in2;
   input [7:0] in1;
   output [31:0] out1;
   input clk;
wire csa_tree_add_39_2_groupi_n_0, csa_tree_add_39_2_groupi_n_1,
     csa_tree_add_39_2_groupi_n_2, csa_tree_add_39_2_groupi_n_3,
     csa_tree_add_39_2_groupi_n_4, csa_tree_add_39_2_groupi_n_5,
     csa_tree_add_39_2_groupi_n_6, csa_tree_add_39_2_groupi_n_7,
     csa_tree_add_39_2_groupi_n_8, csa_tree_add_39_2_groupi_n_9,
     csa_tree_add_39_2_groupi_n_10, csa_tree_add_39_2_groupi_n_12,
     csa_tree_add_39_2_groupi_n_14, csa_tree_add_39_2_groupi_n_15,
     csa_tree_add_39_2_groupi_n_16, csa_tree_add_39_2_groupi_n_17,
     csa_tree_add_39_2_groupi_n_18, csa_tree_add_39_2_groupi_n_19,
     csa_tree_add_39_2_groupi_n_20, csa_tree_add_39_2_groupi_n_21,
     csa_tree_add_39_2_groupi_n_22, csa_tree_add_39_2_groupi_n_23,
     csa_tree_add_39_2_groupi_n_24, csa_tree_add_39_2_groupi_n_25,
     csa_tree_add_39_2_groupi_n_26, csa_tree_add_39_2_groupi_n_27,
     csa_tree_add_39_2_groupi_n_28, csa_tree_add_39_2_groupi_n_29,
     csa_tree_add_39_2_groupi_n_30, csa_tree_add_39_2_groupi_n_31,
     csa_tree_add_39_2_groupi_n_32, csa_tree_add_39_2_groupi_n_33,
     csa_tree_add_39_2_groupi_n_34, csa_tree_add_39_2_groupi_n_35,
     csa_tree_add_39_2_groupi_n_36, csa_tree_add_39_2_groupi_n_37,
     csa_tree_add_39_2_groupi_n_38, csa_tree_add_39_2_groupi_n_39,
     csa_tree_add_39_2_groupi_n_40, csa_tree_add_39_2_groupi_n_41,
     csa_tree_add_39_2_groupi_n_42, csa_tree_add_39_2_groupi_n_43,
     csa_tree_add_39_2_groupi_n_44, csa_tree_add_39_2_groupi_n_45,
     csa_tree_add_39_2_groupi_n_46, csa_tree_add_39_2_groupi_n_47,
     csa_tree_add_39_2_groupi_n_48, csa_tree_add_39_2_groupi_n_49,
     csa_tree_add_39_2_groupi_n_50, csa_tree_add_39_2_groupi_n_51,
     csa_tree_add_39_2_groupi_n_52, csa_tree_add_39_2_groupi_n_53,
     csa_tree_add_39_2_groupi_n_54, csa_tree_add_39_2_groupi_n_55,
     csa_tree_add_39_2_groupi_n_56, csa_tree_add_39_2_groupi_n_57,
     csa_tree_add_39_2_groupi_n_58, csa_tree_add_39_2_groupi_n_59,
     csa_tree_add_39_2_groupi_n_60, csa_tree_add_39_2_groupi_n_61,
     csa_tree_add_39_2_groupi_n_62, csa_tree_add_39_2_groupi_n_63,
     csa_tree_add_39_2_groupi_n_64, csa_tree_add_39_2_groupi_n_65,
     csa_tree_add_39_2_groupi_n_66, csa_tree_add_39_2_groupi_n_67,
     csa_tree_add_39_2_groupi_n_68, csa_tree_add_39_2_groupi_n_69,
     csa_tree_add_39_2_groupi_n_70, csa_tree_add_39_2_groupi_n_71,
     csa_tree_add_39_2_groupi_n_72, csa_tree_add_39_2_groupi_n_73,
     csa_tree_add_39_2_groupi_n_74, csa_tree_add_39_2_groupi_n_75,
     csa_tree_add_39_2_groupi_n_76, csa_tree_add_39_2_groupi_n_77,
     csa_tree_add_39_2_groupi_n_78, csa_tree_add_39_2_groupi_n_79,
     csa_tree_add_39_2_groupi_n_80, csa_tree_add_39_2_groupi_n_81,
     csa_tree_add_39_2_groupi_n_82, csa_tree_add_39_2_groupi_n_83,
     csa_tree_add_39_2_groupi_n_84, csa_tree_add_39_2_groupi_n_85,
     csa_tree_add_39_2_groupi_n_86, csa_tree_add_39_2_groupi_n_87,
     csa_tree_add_39_2_groupi_n_88, csa_tree_add_39_2_groupi_n_89,
     csa_tree_add_39_2_groupi_n_90, csa_tree_add_39_2_groupi_n_91,
     csa_tree_add_39_2_groupi_n_92, csa_tree_add_39_2_groupi_n_93,
     csa_tree_add_39_2_groupi_n_94, csa_tree_add_39_2_groupi_n_95,
     csa_tree_add_39_2_groupi_n_96, csa_tree_add_39_2_groupi_n_97,
     csa_tree_add_39_2_groupi_n_98, csa_tree_add_39_2_groupi_n_99,
     csa_tree_add_39_2_groupi_n_100, csa_tree_add_39_2_groupi_n_101,
     csa_tree_add_39_2_groupi_n_102, csa_tree_add_39_2_groupi_n_105,
     csa_tree_add_39_2_groupi_n_106, csa_tree_add_39_2_groupi_n_107,
     csa_tree_add_39_2_groupi_n_110, csa_tree_add_39_2_groupi_n_111,
     csa_tree_add_39_2_groupi_n_112, csa_tree_add_39_2_groupi_n_117,
     csa_tree_add_39_2_groupi_n_119, csa_tree_add_39_2_groupi_n_120,
     csa_tree_add_39_2_groupi_n_121, csa_tree_add_39_2_groupi_n_122,
     csa_tree_add_39_2_groupi_n_125, csa_tree_add_39_2_groupi_n_126,
     csa_tree_add_39_2_groupi_n_129, csa_tree_add_39_2_groupi_n_130,
     csa_tree_add_39_2_groupi_n_132, csa_tree_add_39_2_groupi_n_134,
     csa_tree_add_39_2_groupi_n_135, csa_tree_add_39_2_groupi_n_137,
     csa_tree_add_39_2_groupi_n_138, csa_tree_add_39_2_groupi_n_139,
     csa_tree_add_39_2_groupi_n_140, csa_tree_add_39_2_groupi_n_141,
     csa_tree_add_39_2_groupi_n_143, csa_tree_add_39_2_groupi_n_144,
     csa_tree_add_39_2_groupi_n_145, csa_tree_add_39_2_groupi_n_148,
     csa_tree_add_39_2_groupi_n_151, csa_tree_add_39_2_groupi_n_152,
     csa_tree_add_39_2_groupi_n_154, csa_tree_add_39_2_groupi_n_155,
     csa_tree_add_39_2_groupi_n_156, csa_tree_add_39_2_groupi_n_157,
     csa_tree_add_39_2_groupi_n_158, csa_tree_add_39_2_groupi_n_159,
     csa_tree_add_39_2_groupi_n_160, csa_tree_add_39_2_groupi_n_161,
     csa_tree_add_39_2_groupi_n_162, csa_tree_add_39_2_groupi_n_163,
     csa_tree_add_39_2_groupi_n_164, csa_tree_add_39_2_groupi_n_165,
     csa_tree_add_39_2_groupi_n_166, csa_tree_add_39_2_groupi_n_167,
     csa_tree_add_39_2_groupi_n_168, csa_tree_add_39_2_groupi_n_169,
     csa_tree_add_39_2_groupi_n_170, csa_tree_add_39_2_groupi_n_171,
     csa_tree_add_39_2_groupi_n_172, csa_tree_add_39_2_groupi_n_173,
     csa_tree_add_39_2_groupi_n_174, csa_tree_add_39_2_groupi_n_175,
     csa_tree_add_39_2_groupi_n_176, csa_tree_add_39_2_groupi_n_177,
     csa_tree_add_39_2_groupi_n_178, csa_tree_add_39_2_groupi_n_179,
     csa_tree_add_39_2_groupi_n_180, csa_tree_add_39_2_groupi_n_181,
     csa_tree_add_39_2_groupi_n_182, csa_tree_add_39_2_groupi_n_183,
     csa_tree_add_39_2_groupi_n_184, csa_tree_add_39_2_groupi_n_185,
     csa_tree_add_39_2_groupi_n_186, csa_tree_add_39_2_groupi_n_190,
     csa_tree_add_39_2_groupi_n_191, csa_tree_add_39_2_groupi_n_192,
     csa_tree_add_39_2_groupi_n_193, csa_tree_add_39_2_groupi_n_194,
     csa_tree_add_39_2_groupi_n_195, csa_tree_add_39_2_groupi_n_196,
     csa_tree_add_39_2_groupi_n_197, csa_tree_add_39_2_groupi_n_198,
     csa_tree_add_39_2_groupi_n_199, csa_tree_add_39_2_groupi_n_200,
     csa_tree_add_39_2_groupi_n_201, csa_tree_add_39_2_groupi_n_202,
     csa_tree_add_39_2_groupi_n_203, csa_tree_add_39_2_groupi_n_208,
     csa_tree_add_39_2_groupi_n_213, csa_tree_add_39_2_groupi_n_214,
     csa_tree_add_39_2_groupi_n_215, csa_tree_add_39_2_groupi_n_216,
     csa_tree_add_39_2_groupi_n_217, csa_tree_add_39_2_groupi_n_218,
     csa_tree_add_39_2_groupi_n_221, csa_tree_add_39_2_groupi_n_222,
     csa_tree_add_39_2_groupi_n_224, csa_tree_add_39_2_groupi_n_225,
     csa_tree_add_39_2_groupi_n_226, csa_tree_add_39_2_groupi_n_227,
     csa_tree_add_39_2_groupi_n_228, csa_tree_add_39_2_groupi_n_229,
     csa_tree_add_39_2_groupi_n_230, csa_tree_add_39_2_groupi_n_231,
     csa_tree_add_39_2_groupi_n_232, csa_tree_add_39_2_groupi_n_233,
     csa_tree_add_39_2_groupi_n_234, csa_tree_add_39_2_groupi_n_239,
     csa_tree_add_39_2_groupi_n_240, csa_tree_add_39_2_groupi_n_241,
     csa_tree_add_39_2_groupi_n_242, csa_tree_add_39_2_groupi_n_245,
     csa_tree_add_39_2_groupi_n_247, csa_tree_add_39_2_groupi_n_249,
     csa_tree_add_39_2_groupi_n_250, csa_tree_add_39_2_groupi_n_251,
     csa_tree_add_39_2_groupi_n_252, csa_tree_add_39_2_groupi_n_253,
     csa_tree_add_39_2_groupi_n_256, csa_tree_add_39_2_groupi_n_257,
     csa_tree_add_39_2_groupi_n_258, csa_tree_add_39_2_groupi_n_259,
     csa_tree_add_39_2_groupi_n_262, csa_tree_add_39_2_groupi_n_263,
     csa_tree_add_39_2_groupi_n_265, csa_tree_add_39_2_groupi_n_266,
     csa_tree_add_39_2_groupi_n_267, csa_tree_add_39_2_groupi_n_268,
     csa_tree_add_39_2_groupi_n_269, csa_tree_add_39_2_groupi_n_272,
     csa_tree_add_39_2_groupi_n_273, csa_tree_add_39_2_groupi_n_274,
     csa_tree_add_39_2_groupi_n_275, csa_tree_add_39_2_groupi_n_278,
     csa_tree_add_39_2_groupi_n_279, csa_tree_add_39_2_groupi_n_280,
     csa_tree_add_39_2_groupi_n_281, csa_tree_add_39_2_groupi_n_301,
     csa_tree_add_39_2_groupi_n_302, csa_tree_add_39_2_groupi_n_304,
     csa_tree_add_39_2_groupi_n_306, csa_tree_add_39_2_groupi_n_308,
     csa_tree_add_39_2_groupi_n_310, csa_tree_add_39_2_groupi_n_312,
     csa_tree_add_39_2_groupi_n_314, csa_tree_add_39_2_groupi_n_316,
     csa_tree_add_39_2_groupi_n_318, n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8,
     n_9, n_10, n_11, n_12, n_13, clk, n_47, n_48, n_49, n_50, n_51, n_52, n_53,
     n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64, n_65,
     n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76, n_77,
     n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_102, n_103, n_104, n_105,
     n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116;
 reg out1_6_L0_reg_N30;
 always @(posedge clk)
         out1_6_L0_reg_N30 <= n_8;
 assign {out1[25]} = out1_6_L0_reg_N30;
 reg out1_7_L0_reg_N30;
 always @(posedge clk)
         out1_7_L0_reg_N30 <= n_9;
 assign {out1[24]} = out1_7_L0_reg_N30;
 reg out1_8_L0_reg_N30;
 always @(posedge clk)
         out1_8_L0_reg_N30 <= n_12;
 assign {out1[23]} = out1_8_L0_reg_N30;
 reg out1_9_L0_reg_N30;
 always @(posedge clk)
         out1_9_L0_reg_N30 <= n_5;
 assign {out1[22]} = out1_9_L0_reg_N30;
 reg out1_10_L0_reg_N30;
 always @(posedge clk)
         out1_10_L0_reg_N30 <= n_6;
 assign {out1[21]} = out1_10_L0_reg_N30;
 reg out1_11_L0_reg_N30;
 always @(posedge clk)
         out1_11_L0_reg_N30 <= n_3;
 assign {out1[20]} = out1_11_L0_reg_N30;
 reg out1_12_L0_reg_N30;
 always @(posedge clk)
         out1_12_L0_reg_N30 <= n_4;
 assign {out1[19]} = out1_12_L0_reg_N30;
 reg out1_13_L0_reg_N30;
 always @(posedge clk)
         out1_13_L0_reg_N30 <= n_7;
 assign {out1[18]} = out1_13_L0_reg_N30;
 reg out1_14_L0_reg_N30;
 always @(posedge clk)
         out1_14_L0_reg_N30 <= n_10;
 assign {out1[17]} = out1_14_L0_reg_N30;
 reg out1_15_L0_reg_N30;
 always @(posedge clk)
         if ({in3[16]})
         out1_15_L0_reg_N30 <= n_54;
     else
         out1_15_L0_reg_N30 <= csa_tree_add_39_2_groupi_n_301;
 assign {out1[16]} = out1_15_L0_reg_N30;
 reg out1_16_L0_reg_N30;
 always @(posedge clk)
         out1_16_L0_reg_N30 <= n_55;
 assign {out1[15]} = out1_16_L0_reg_N30;
 reg out1_17_L0_reg_N30;
 always @(posedge clk)
         out1_17_L0_reg_N30 <= n_56;
 assign {out1[14]} = out1_17_L0_reg_N30;
 reg out1_18_L0_reg_N30;
 always @(posedge clk)
         out1_18_L0_reg_N30 <= n_58;
 assign {out1[13]} = out1_18_L0_reg_N30;
 reg out1_19_L0_reg_N30;
 always @(posedge clk)
         out1_19_L0_reg_N30 <= n_60;
 assign {out1[12]} = out1_19_L0_reg_N30;
 reg out1_20_L0_reg_N30;
 always @(posedge clk)
         out1_20_L0_reg_N30 <= n_62;
 assign {out1[11]} = out1_20_L0_reg_N30;
 reg out1_21_L0_reg_N30;
 always @(posedge clk)
         out1_21_L0_reg_N30 <= n_64;
 assign {out1[10]} = out1_21_L0_reg_N30;
 reg out1_22_L0_reg_N30;
 always @(posedge clk)
         out1_22_L0_reg_N30 <= n_66;
 assign {out1[9]} = out1_22_L0_reg_N30;
 reg out1_23_L0_reg_N30;
 always @(posedge clk)
         out1_23_L0_reg_N30 <= n_68;
 assign {out1[8]} = out1_23_L0_reg_N30;
 reg out1_24_L0_reg_N30;
 always @(posedge clk)
         out1_24_L0_reg_N30 <= n_70;
 assign {out1[7]} = out1_24_L0_reg_N30;
 reg out1_25_L0_reg_N30;
 always @(posedge clk)
         out1_25_L0_reg_N30 <= n_72;
 assign {out1[6]} = out1_25_L0_reg_N30;
 reg out1_26_L0_reg_N30;
 always @(posedge clk)
         out1_26_L0_reg_N30 <= n_74;
 assign {out1[5]} = out1_26_L0_reg_N30;
 reg out1_27_L0_reg_N30;
 always @(posedge clk)
         out1_27_L0_reg_N30 <= n_76;
 assign {out1[4]} = out1_27_L0_reg_N30;
 reg out1_28_L0_reg_N30;
 always @(posedge clk)
         out1_28_L0_reg_N30 <= n_78;
 assign {out1[3]} = out1_28_L0_reg_N30;
 reg out1_29_L0_reg_N30;
 always @(posedge clk)
         out1_29_L0_reg_N30 <= n_83;
 assign {out1[2]} = out1_29_L0_reg_N30;
 reg out1_30_L0_reg_N30;
 always @(posedge clk)
         out1_30_L0_reg_N30 <= n_1;
 assign {out1[1]} = out1_30_L0_reg_N30;
 reg out1_31_L0_reg_N30;
 always @(posedge clk)
         out1_31_L0_reg_N30 <= n_11;
 assign {out1[0]} = out1_31_L0_reg_N30;
 reg retime_s1_1_reg_reg_N30;
 always @(posedge clk)
         retime_s1_1_reg_reg_N30 <= {in3[30]};
 assign n_47 = retime_s1_1_reg_reg_N30;
 reg retime_s1_2_reg_reg_N30;
 always @(posedge clk)
         retime_s1_2_reg_reg_N30 <= {in3[31]};
 assign n_48 = retime_s1_2_reg_reg_N30;
 reg retime_s1_3_reg_reg_N30;
 always @(posedge clk)
         retime_s1_3_reg_reg_N30 <= {in3[28]};
 assign n_49 = retime_s1_3_reg_reg_N30;
 reg retime_s1_4_reg_reg_N30;
 always @(posedge clk)
         retime_s1_4_reg_reg_N30 <= {in3[29]};
 assign n_50 = retime_s1_4_reg_reg_N30;
 reg retime_s1_5_reg_reg_N30;
 always @(posedge clk)
         retime_s1_5_reg_reg_N30 <= {in3[27]};
 assign n_51 = retime_s1_5_reg_reg_N30;
 reg retime_s1_6_reg_reg_N30;
 always @(posedge clk)
         retime_s1_6_reg_reg_N30 <= {in3[26]};
 assign n_52 = retime_s1_6_reg_reg_N30;
 reg retime_s1_7_reg_reg_N30;
 always @(posedge clk)
         retime_s1_7_reg_reg_N30 <= n_13;
 assign n_53 = retime_s1_7_reg_reg_N30;
 assign csa_tree_add_39_2_groupi_n_20 = ({in2[3]} & {in1[1]});
 assign csa_tree_add_39_2_groupi_n_318 = ~({in3[24]} & ~csa_tree_add_39_2_groupi_n_316);
 assign csa_tree_add_39_2_groupi_n_316 = ~({in3[23]} & ~csa_tree_add_39_2_groupi_n_314);
 assign csa_tree_add_39_2_groupi_n_314 = ~({in3[22]} & ~csa_tree_add_39_2_groupi_n_312);
 assign csa_tree_add_39_2_groupi_n_312 = ~({in3[21]} & ~csa_tree_add_39_2_groupi_n_310);
 assign csa_tree_add_39_2_groupi_n_310 = ~({in3[20]} & ~csa_tree_add_39_2_groupi_n_308);
 assign csa_tree_add_39_2_groupi_n_308 = ~({in3[19]} & ~csa_tree_add_39_2_groupi_n_306);
 assign csa_tree_add_39_2_groupi_n_306 = ~({in3[18]} & ~csa_tree_add_39_2_groupi_n_304);
 assign csa_tree_add_39_2_groupi_n_304 = ~({in3[17]} & ~csa_tree_add_39_2_groupi_n_302);
 assign csa_tree_add_39_2_groupi_n_302 = ~(csa_tree_add_39_2_groupi_n_301 & {in3[16]});
 assign csa_tree_add_39_2_groupi_n_280 = ((csa_tree_add_39_2_groupi_n_256 & csa_tree_add_39_2_groupi_n_259)
    | ((csa_tree_add_39_2_groupi_n_259 & csa_tree_add_39_2_groupi_n_234) | (csa_tree_add_39_2_groupi_n_234
    & csa_tree_add_39_2_groupi_n_256)));
 assign csa_tree_add_39_2_groupi_n_281 = (csa_tree_add_39_2_groupi_n_259 ^ (csa_tree_add_39_2_groupi_n_234
    ^ csa_tree_add_39_2_groupi_n_256));
 assign csa_tree_add_39_2_groupi_n_278 = ((csa_tree_add_39_2_groupi_n_258 & csa_tree_add_39_2_groupi_n_263)
    | ((csa_tree_add_39_2_groupi_n_263 & csa_tree_add_39_2_groupi_n_242) | (csa_tree_add_39_2_groupi_n_242
    & csa_tree_add_39_2_groupi_n_258)));
 assign csa_tree_add_39_2_groupi_n_279 = (csa_tree_add_39_2_groupi_n_263 ^ (csa_tree_add_39_2_groupi_n_242
    ^ csa_tree_add_39_2_groupi_n_258));
 assign csa_tree_add_39_2_groupi_n_274 = ((csa_tree_add_39_2_groupi_n_249 & csa_tree_add_39_2_groupi_n_257)
    | ((csa_tree_add_39_2_groupi_n_257 & csa_tree_add_39_2_groupi_n_232) | (csa_tree_add_39_2_groupi_n_232
    & csa_tree_add_39_2_groupi_n_249)));
 assign csa_tree_add_39_2_groupi_n_275 = (csa_tree_add_39_2_groupi_n_257 ^ (csa_tree_add_39_2_groupi_n_232
    ^ csa_tree_add_39_2_groupi_n_249));
 assign csa_tree_add_39_2_groupi_n_272 = ((csa_tree_add_39_2_groupi_n_250 & csa_tree_add_39_2_groupi_n_225)
    | ((csa_tree_add_39_2_groupi_n_225 & csa_tree_add_39_2_groupi_n_240) | (csa_tree_add_39_2_groupi_n_240
    & csa_tree_add_39_2_groupi_n_250)));
 assign csa_tree_add_39_2_groupi_n_273 = (csa_tree_add_39_2_groupi_n_225 ^ (csa_tree_add_39_2_groupi_n_240
    ^ csa_tree_add_39_2_groupi_n_250));
 assign csa_tree_add_39_2_groupi_n_268 = ((csa_tree_add_39_2_groupi_n_262 & csa_tree_add_39_2_groupi_n_241)
    | ((csa_tree_add_39_2_groupi_n_241 & csa_tree_add_39_2_groupi_n_229) | (csa_tree_add_39_2_groupi_n_229
    & csa_tree_add_39_2_groupi_n_262)));
 assign csa_tree_add_39_2_groupi_n_269 = (csa_tree_add_39_2_groupi_n_241 ^ (csa_tree_add_39_2_groupi_n_229
    ^ csa_tree_add_39_2_groupi_n_262));
 assign csa_tree_add_39_2_groupi_n_266 = ((csa_tree_add_39_2_groupi_n_228 & csa_tree_add_39_2_groupi_n_197)
    | ((csa_tree_add_39_2_groupi_n_197 & csa_tree_add_39_2_groupi_n_227) | (csa_tree_add_39_2_groupi_n_227
    & csa_tree_add_39_2_groupi_n_228)));
 assign csa_tree_add_39_2_groupi_n_267 = (csa_tree_add_39_2_groupi_n_197 ^ (csa_tree_add_39_2_groupi_n_227
    ^ csa_tree_add_39_2_groupi_n_228));
 assign csa_tree_add_39_2_groupi_n_265 = ~(csa_tree_add_39_2_groupi_n_253 & ~(csa_tree_add_39_2_groupi_n_218
    & csa_tree_add_39_2_groupi_n_230));
 assign csa_tree_add_39_2_groupi_n_262 = ((csa_tree_add_39_2_groupi_n_233 & csa_tree_add_39_2_groupi_n_162)
    | ((csa_tree_add_39_2_groupi_n_162 & csa_tree_add_39_2_groupi_n_215) | (csa_tree_add_39_2_groupi_n_215
    & csa_tree_add_39_2_groupi_n_233)));
 assign csa_tree_add_39_2_groupi_n_263 = (csa_tree_add_39_2_groupi_n_162 ^ (csa_tree_add_39_2_groupi_n_215
    ^ csa_tree_add_39_2_groupi_n_233));
 assign csa_tree_add_39_2_groupi_n_258 = ((csa_tree_add_39_2_groupi_n_231 & csa_tree_add_39_2_groupi_n_213)
    | ((csa_tree_add_39_2_groupi_n_213 & csa_tree_add_39_2_groupi_n_216) | (csa_tree_add_39_2_groupi_n_216
    & csa_tree_add_39_2_groupi_n_231)));
 assign csa_tree_add_39_2_groupi_n_259 = (csa_tree_add_39_2_groupi_n_213 ^ (csa_tree_add_39_2_groupi_n_216
    ^ csa_tree_add_39_2_groupi_n_231));
 assign csa_tree_add_39_2_groupi_n_256 = ((csa_tree_add_39_2_groupi_n_239 & csa_tree_add_39_2_groupi_n_193)
    | ((csa_tree_add_39_2_groupi_n_193 & csa_tree_add_39_2_groupi_n_214) | (csa_tree_add_39_2_groupi_n_214
    & csa_tree_add_39_2_groupi_n_239)));
 assign csa_tree_add_39_2_groupi_n_257 = (csa_tree_add_39_2_groupi_n_193 ^ (csa_tree_add_39_2_groupi_n_214
    ^ csa_tree_add_39_2_groupi_n_239));
 assign csa_tree_add_39_2_groupi_n_253 = ~(csa_tree_add_39_2_groupi_n_245 & (csa_tree_add_39_2_groupi_n_218
    | csa_tree_add_39_2_groupi_n_230));
 assign csa_tree_add_39_2_groupi_n_251 = ((csa_tree_add_39_2_groupi_n_226 & csa_tree_add_39_2_groupi_n_157)
    | ((csa_tree_add_39_2_groupi_n_157 & csa_tree_add_39_2_groupi_n_160) | (csa_tree_add_39_2_groupi_n_160
    & csa_tree_add_39_2_groupi_n_226)));
 assign csa_tree_add_39_2_groupi_n_252 = (csa_tree_add_39_2_groupi_n_157 ^ (csa_tree_add_39_2_groupi_n_160
    ^ csa_tree_add_39_2_groupi_n_226));
 assign csa_tree_add_39_2_groupi_n_249 = ((csa_tree_add_39_2_groupi_n_217 & csa_tree_add_39_2_groupi_n_194)
    | ((csa_tree_add_39_2_groupi_n_194 & csa_tree_add_39_2_groupi_n_181) | (csa_tree_add_39_2_groupi_n_181
    & csa_tree_add_39_2_groupi_n_217)));
 assign csa_tree_add_39_2_groupi_n_250 = (csa_tree_add_39_2_groupi_n_194 ^ (csa_tree_add_39_2_groupi_n_181
    ^ csa_tree_add_39_2_groupi_n_217));
 assign csa_tree_add_39_2_groupi_n_247 = ~(csa_tree_add_39_2_groupi_n_17 & ~(csa_tree_add_39_2_groupi_n_185
    & csa_tree_add_39_2_groupi_n_200));
 assign csa_tree_add_39_2_groupi_n_245 = ~csa_tree_add_39_2_groupi_n_16;
 assign csa_tree_add_39_2_groupi_n_241 = ((csa_tree_add_39_2_groupi_n_156 & csa_tree_add_39_2_groupi_n_178)
    | ((csa_tree_add_39_2_groupi_n_178 & csa_tree_add_39_2_groupi_n_174) | (csa_tree_add_39_2_groupi_n_174
    & csa_tree_add_39_2_groupi_n_156)));
 assign csa_tree_add_39_2_groupi_n_242 = (csa_tree_add_39_2_groupi_n_178 ^ (csa_tree_add_39_2_groupi_n_174
    ^ csa_tree_add_39_2_groupi_n_156));
 assign csa_tree_add_39_2_groupi_n_239 = ((csa_tree_add_39_2_groupi_n_177 & csa_tree_add_39_2_groupi_n_151)
    | ((csa_tree_add_39_2_groupi_n_151 & csa_tree_add_39_2_groupi_n_173) | (csa_tree_add_39_2_groupi_n_173
    & csa_tree_add_39_2_groupi_n_177)));
 assign csa_tree_add_39_2_groupi_n_240 = (csa_tree_add_39_2_groupi_n_151 ^ (csa_tree_add_39_2_groupi_n_173
    ^ csa_tree_add_39_2_groupi_n_177));
 assign csa_tree_add_39_2_groupi_n_233 = ((csa_tree_add_39_2_groupi_n_175 & csa_tree_add_39_2_groupi_n_163)
    | ((csa_tree_add_39_2_groupi_n_163 & csa_tree_add_39_2_groupi_n_179) | (csa_tree_add_39_2_groupi_n_179
    & csa_tree_add_39_2_groupi_n_175)));
 assign csa_tree_add_39_2_groupi_n_234 = (csa_tree_add_39_2_groupi_n_163 ^ (csa_tree_add_39_2_groupi_n_179
    ^ csa_tree_add_39_2_groupi_n_175));
 assign csa_tree_add_39_2_groupi_n_231 = ((csa_tree_add_39_2_groupi_n_164 & csa_tree_add_39_2_groupi_n_176)
    | ((csa_tree_add_39_2_groupi_n_176 & csa_tree_add_39_2_groupi_n_172) | (csa_tree_add_39_2_groupi_n_172
    & csa_tree_add_39_2_groupi_n_164)));
 assign csa_tree_add_39_2_groupi_n_232 = (csa_tree_add_39_2_groupi_n_176 ^ (csa_tree_add_39_2_groupi_n_172
    ^ csa_tree_add_39_2_groupi_n_164));
 assign csa_tree_add_39_2_groupi_n_230 = ~csa_tree_add_39_2_groupi_n_222;
 assign csa_tree_add_39_2_groupi_n_228 = ((csa_tree_add_39_2_groupi_n_198 & csa_tree_add_39_2_groupi_n_155)
    | ((csa_tree_add_39_2_groupi_n_155 & csa_tree_add_39_2_groupi_n_166) | (csa_tree_add_39_2_groupi_n_166
    & csa_tree_add_39_2_groupi_n_198)));
 assign csa_tree_add_39_2_groupi_n_229 = (csa_tree_add_39_2_groupi_n_155 ^ (csa_tree_add_39_2_groupi_n_166
    ^ csa_tree_add_39_2_groupi_n_198));
 assign csa_tree_add_39_2_groupi_n_226 = ((csa_tree_add_39_2_groupi_n_158 & csa_tree_add_39_2_groupi_n_79)
    | ((csa_tree_add_39_2_groupi_n_79 & csa_tree_add_39_2_groupi_n_165) | (csa_tree_add_39_2_groupi_n_165
    & csa_tree_add_39_2_groupi_n_158)));
 assign csa_tree_add_39_2_groupi_n_227 = (csa_tree_add_39_2_groupi_n_79 ^ (csa_tree_add_39_2_groupi_n_165
    ^ csa_tree_add_39_2_groupi_n_158));
 assign csa_tree_add_39_2_groupi_n_225 = ~(csa_tree_add_39_2_groupi_n_224 & csa_tree_add_39_2_groupi_n_186);
 assign csa_tree_add_39_2_groupi_n_224 = ~(csa_tree_add_39_2_groupi_n_15 & csa_tree_add_39_2_groupi_n_184);
 assign csa_tree_add_39_2_groupi_n_222 = ~(csa_tree_add_39_2_groupi_n_203 | csa_tree_add_39_2_groupi_n_192);
 assign csa_tree_add_39_2_groupi_n_221 = ~(csa_tree_add_39_2_groupi_n_168 & (csa_tree_add_39_2_groupi_n_202
    | csa_tree_add_39_2_groupi_n_170));
 assign csa_tree_add_39_2_groupi_n_217 = ((csa_tree_add_39_2_groupi_n_152 & csa_tree_add_39_2_groupi_n_0)
    | ((csa_tree_add_39_2_groupi_n_0 & csa_tree_add_39_2_groupi_n_139) | (csa_tree_add_39_2_groupi_n_139
    & csa_tree_add_39_2_groupi_n_152)));
 assign csa_tree_add_39_2_groupi_n_218 = (csa_tree_add_39_2_groupi_n_0 ^ (csa_tree_add_39_2_groupi_n_139
    ^ csa_tree_add_39_2_groupi_n_152));
 assign csa_tree_add_39_2_groupi_n_215 = ((csa_tree_add_39_2_groupi_n_171 & csa_tree_add_39_2_groupi_n_81)
    | ((csa_tree_add_39_2_groupi_n_81 & csa_tree_add_39_2_groupi_n_101) | (csa_tree_add_39_2_groupi_n_101
    & csa_tree_add_39_2_groupi_n_171)));
 assign csa_tree_add_39_2_groupi_n_216 = (csa_tree_add_39_2_groupi_n_81 ^ (csa_tree_add_39_2_groupi_n_101
    ^ csa_tree_add_39_2_groupi_n_171));
 assign csa_tree_add_39_2_groupi_n_213 = ((csa_tree_add_39_2_groupi_n_180 & csa_tree_add_39_2_groupi_n_110)
    | ((csa_tree_add_39_2_groupi_n_110 & n_112) | (n_112 & csa_tree_add_39_2_groupi_n_180)));
 assign csa_tree_add_39_2_groupi_n_214 = (csa_tree_add_39_2_groupi_n_110 ^ (n_112 ^ csa_tree_add_39_2_groupi_n_180));
 assign csa_tree_add_39_2_groupi_n_208 = (csa_tree_add_39_2_groupi_n_185 | csa_tree_add_39_2_groupi_n_200);
 assign csa_tree_add_39_2_groupi_n_203 = ~(csa_tree_add_39_2_groupi_n_7 | csa_tree_add_39_2_groupi_n_169);
 assign csa_tree_add_39_2_groupi_n_200 = ~csa_tree_add_39_2_groupi_n_201;
 assign csa_tree_add_39_2_groupi_n_197 = ((csa_tree_add_39_2_groupi_n_161 & csa_tree_add_39_2_groupi_n_46)
    | ((csa_tree_add_39_2_groupi_n_46 & csa_tree_add_39_2_groupi_n_82) | (csa_tree_add_39_2_groupi_n_82 &
    csa_tree_add_39_2_groupi_n_161)));
 assign csa_tree_add_39_2_groupi_n_198 = (csa_tree_add_39_2_groupi_n_46 ^ (csa_tree_add_39_2_groupi_n_82
    ^ csa_tree_add_39_2_groupi_n_161));
 assign csa_tree_add_39_2_groupi_n_195 = ((csa_tree_add_39_2_groupi_n_159 & csa_tree_add_39_2_groupi_n_45)
    | ((csa_tree_add_39_2_groupi_n_45 & {in3[14]}) | ({in3[14]} & csa_tree_add_39_2_groupi_n_159)));
 assign csa_tree_add_39_2_groupi_n_196 = (csa_tree_add_39_2_groupi_n_45 ^ ({in3[14]} ^ csa_tree_add_39_2_groupi_n_159));
 assign csa_tree_add_39_2_groupi_n_201 = ((csa_tree_add_39_2_groupi_n_129 & csa_tree_add_39_2_groupi_n_42)
    | ((csa_tree_add_39_2_groupi_n_42 & csa_tree_add_39_2_groupi_n_112) | (csa_tree_add_39_2_groupi_n_112
    & csa_tree_add_39_2_groupi_n_129)));
 assign csa_tree_add_39_2_groupi_n_202 = (csa_tree_add_39_2_groupi_n_42 ^ (csa_tree_add_39_2_groupi_n_112
    ^ csa_tree_add_39_2_groupi_n_129));
 assign csa_tree_add_39_2_groupi_n_193 = ((csa_tree_add_39_2_groupi_n_122 & csa_tree_add_39_2_groupi_n_84)
    | ((csa_tree_add_39_2_groupi_n_84 & csa_tree_add_39_2_groupi_n_138) | (csa_tree_add_39_2_groupi_n_138
    & csa_tree_add_39_2_groupi_n_122)));
 assign csa_tree_add_39_2_groupi_n_194 = (csa_tree_add_39_2_groupi_n_84 ^ (csa_tree_add_39_2_groupi_n_138
    ^ csa_tree_add_39_2_groupi_n_122));
 assign csa_tree_add_39_2_groupi_n_192 = (csa_tree_add_39_2_groupi_n_135 & n_113);
 assign csa_tree_add_39_2_groupi_n_199 = (csa_tree_add_39_2_groupi_n_135 ^ n_113);
 assign csa_tree_add_39_2_groupi_n_191 = ~((csa_tree_add_39_2_groupi_n_183 & ~csa_tree_add_39_2_groupi_n_182)
    | (n_109 & csa_tree_add_39_2_groupi_n_182));
 assign csa_tree_add_39_2_groupi_n_190 = ~(csa_tree_add_39_2_groupi_n_145 & (n_111 | csa_tree_add_39_2_groupi_n_148));
 assign csa_tree_add_39_2_groupi_n_186 = ~(csa_tree_add_39_2_groupi_n_182 & csa_tree_add_39_2_groupi_n_183);
 assign csa_tree_add_39_2_groupi_n_183 = ~n_109;
 assign csa_tree_add_39_2_groupi_n_180 = ((csa_tree_add_39_2_groupi_n_2 & csa_tree_add_39_2_groupi_n_83)
    | ((csa_tree_add_39_2_groupi_n_83 & csa_tree_add_39_2_groupi_n_77) | (csa_tree_add_39_2_groupi_n_77 &
    csa_tree_add_39_2_groupi_n_2)));
 assign csa_tree_add_39_2_groupi_n_181 = (csa_tree_add_39_2_groupi_n_83 ^ (csa_tree_add_39_2_groupi_n_77
    ^ csa_tree_add_39_2_groupi_n_2));
 assign csa_tree_add_39_2_groupi_n_178 = ((csa_tree_add_39_2_groupi_n_87 & csa_tree_add_39_2_groupi_n_41)
    | ((csa_tree_add_39_2_groupi_n_41 & {in3[9]}) | ({in3[9]} & csa_tree_add_39_2_groupi_n_87)));
 assign csa_tree_add_39_2_groupi_n_179 = (csa_tree_add_39_2_groupi_n_41 ^ ({in3[9]} ^ csa_tree_add_39_2_groupi_n_87));
 assign csa_tree_add_39_2_groupi_n_176 = ((csa_tree_add_39_2_groupi_n_53 & csa_tree_add_39_2_groupi_n_43)
    | ((csa_tree_add_39_2_groupi_n_43 & csa_tree_add_39_2_groupi_n_71) | (csa_tree_add_39_2_groupi_n_71 &
    csa_tree_add_39_2_groupi_n_53)));
 assign csa_tree_add_39_2_groupi_n_177 = (csa_tree_add_39_2_groupi_n_43 ^ (csa_tree_add_39_2_groupi_n_71
    ^ csa_tree_add_39_2_groupi_n_53));
 assign csa_tree_add_39_2_groupi_n_174 = ((csa_tree_add_39_2_groupi_n_50 & csa_tree_add_39_2_groupi_n_48)
    | ((csa_tree_add_39_2_groupi_n_48 & csa_tree_add_39_2_groupi_n_44) | (csa_tree_add_39_2_groupi_n_44 &
    csa_tree_add_39_2_groupi_n_50)));
 assign csa_tree_add_39_2_groupi_n_175 = (csa_tree_add_39_2_groupi_n_48 ^ (csa_tree_add_39_2_groupi_n_44
    ^ csa_tree_add_39_2_groupi_n_50));
 assign csa_tree_add_39_2_groupi_n_184 = ((csa_tree_add_39_2_groupi_n_102 & csa_tree_add_39_2_groupi_n_19)
    | ((csa_tree_add_39_2_groupi_n_19 & csa_tree_add_39_2_groupi_n_18) | (csa_tree_add_39_2_groupi_n_18 &
    csa_tree_add_39_2_groupi_n_102)));
 assign csa_tree_add_39_2_groupi_n_185 = (csa_tree_add_39_2_groupi_n_19 ^ (csa_tree_add_39_2_groupi_n_18
    ^ csa_tree_add_39_2_groupi_n_102));
 assign csa_tree_add_39_2_groupi_n_173 = ((csa_tree_add_39_2_groupi_n_54 & csa_tree_add_39_2_groupi_n_76)
    | ((csa_tree_add_39_2_groupi_n_76 & csa_tree_add_39_2_groupi_n_47) | (csa_tree_add_39_2_groupi_n_47 &
    csa_tree_add_39_2_groupi_n_54)));
 assign csa_tree_add_39_2_groupi_n_182 = (csa_tree_add_39_2_groupi_n_76 ^ (csa_tree_add_39_2_groupi_n_47
    ^ csa_tree_add_39_2_groupi_n_54));
 assign csa_tree_add_39_2_groupi_n_171 = ((csa_tree_add_39_2_groupi_n_85 & csa_tree_add_39_2_groupi_n_39)
    | ((csa_tree_add_39_2_groupi_n_39 & csa_tree_add_39_2_groupi_n_80) | (csa_tree_add_39_2_groupi_n_80 &
    csa_tree_add_39_2_groupi_n_85)));
 assign csa_tree_add_39_2_groupi_n_172 = (csa_tree_add_39_2_groupi_n_39 ^ (csa_tree_add_39_2_groupi_n_80
    ^ csa_tree_add_39_2_groupi_n_85));
 assign csa_tree_add_39_2_groupi_n_170 = ~(csa_tree_add_39_2_groupi_n_167 | csa_tree_add_39_2_groupi_n_134);
 assign csa_tree_add_39_2_groupi_n_169 = ~(csa_tree_add_39_2_groupi_n_135 | n_113);
 assign csa_tree_add_39_2_groupi_n_168 = ~(csa_tree_add_39_2_groupi_n_167 & csa_tree_add_39_2_groupi_n_134);
 assign csa_tree_add_39_2_groupi_n_167 = ~csa_tree_add_39_2_groupi_n_4;
 assign csa_tree_add_39_2_groupi_n_165 = ((csa_tree_add_39_2_groupi_n_88 & csa_tree_add_39_2_groupi_n_49)
    | ((csa_tree_add_39_2_groupi_n_49 & {in3[11]}) | ({in3[11]} & csa_tree_add_39_2_groupi_n_88)));
 assign csa_tree_add_39_2_groupi_n_166 = (csa_tree_add_39_2_groupi_n_49 ^ ({in3[11]} ^ csa_tree_add_39_2_groupi_n_88));
 assign csa_tree_add_39_2_groupi_n_163 = ((csa_tree_add_39_2_groupi_n_52 & csa_tree_add_39_2_groupi_n_74)
    | ((csa_tree_add_39_2_groupi_n_74 & csa_tree_add_39_2_groupi_n_70) | (csa_tree_add_39_2_groupi_n_70 &
    csa_tree_add_39_2_groupi_n_52)));
 assign csa_tree_add_39_2_groupi_n_164 = (csa_tree_add_39_2_groupi_n_74 ^ (csa_tree_add_39_2_groupi_n_70
    ^ csa_tree_add_39_2_groupi_n_52));
 assign csa_tree_add_39_2_groupi_n_161 = ((csa_tree_add_39_2_groupi_n_51 & csa_tree_add_39_2_groupi_n_40)
    | ((csa_tree_add_39_2_groupi_n_40 & csa_tree_add_39_2_groupi_n_75) | (csa_tree_add_39_2_groupi_n_75 &
    csa_tree_add_39_2_groupi_n_51)));
 assign csa_tree_add_39_2_groupi_n_162 = (csa_tree_add_39_2_groupi_n_40 ^ (csa_tree_add_39_2_groupi_n_75
    ^ csa_tree_add_39_2_groupi_n_51));
 assign csa_tree_add_39_2_groupi_n_159 = ((csa_tree_add_39_2_groupi_n_57 & {in3[13]}) | (({in3[13]} &
    csa_tree_add_39_2_groupi_n_73) | (csa_tree_add_39_2_groupi_n_73 & csa_tree_add_39_2_groupi_n_57)));
 assign csa_tree_add_39_2_groupi_n_160 = ({in3[13]} ^ (csa_tree_add_39_2_groupi_n_73 ^ csa_tree_add_39_2_groupi_n_57));
 assign csa_tree_add_39_2_groupi_n_157 = ((csa_tree_add_39_2_groupi_n_56 & csa_tree_add_39_2_groupi_n_72)
    | ((csa_tree_add_39_2_groupi_n_72 & {in3[12]}) | ({in3[12]} & csa_tree_add_39_2_groupi_n_56)));
 assign csa_tree_add_39_2_groupi_n_158 = (csa_tree_add_39_2_groupi_n_72 ^ ({in3[12]} ^ csa_tree_add_39_2_groupi_n_56));
 assign csa_tree_add_39_2_groupi_n_155 = ((csa_tree_add_39_2_groupi_n_86 & csa_tree_add_39_2_groupi_n_69)
    | ((csa_tree_add_39_2_groupi_n_69 & {in3[10]}) | ({in3[10]} & csa_tree_add_39_2_groupi_n_86)));
 assign csa_tree_add_39_2_groupi_n_156 = (csa_tree_add_39_2_groupi_n_69 ^ ({in3[10]} ^ csa_tree_add_39_2_groupi_n_86));
 assign csa_tree_add_39_2_groupi_n_154 = ~(csa_tree_add_39_2_groupi_n_9 & (csa_tree_add_39_2_groupi_n_125
    | csa_tree_add_39_2_groupi_n_137));
 assign csa_tree_add_39_2_groupi_n_152 = ~(csa_tree_add_39_2_groupi_n_143 & csa_tree_add_39_2_groupi_n_5);
 assign csa_tree_add_39_2_groupi_n_151 = ~(csa_tree_add_39_2_groupi_n_144 & ~csa_tree_add_39_2_groupi_n_117);
 assign csa_tree_add_39_2_groupi_n_148 = ~(csa_tree_add_39_2_groupi_n_141 | csa_tree_add_39_2_groupi_n_1);
 assign csa_tree_add_39_2_groupi_n_145 = ~(csa_tree_add_39_2_groupi_n_141 & csa_tree_add_39_2_groupi_n_1);
 assign csa_tree_add_39_2_groupi_n_144 = ~(csa_tree_add_39_2_groupi_n_65 & ~(csa_tree_add_39_2_groupi_n_90
    & csa_tree_add_39_2_groupi_n_93));
 assign csa_tree_add_39_2_groupi_n_143 = ~(csa_tree_add_39_2_groupi_n_6 & csa_tree_add_39_2_groupi_n_67);
 assign csa_tree_add_39_2_groupi_n_141 = ~csa_tree_add_39_2_groupi_n_132;
 assign csa_tree_add_39_2_groupi_n_138 = (csa_tree_add_39_2_groupi_n_55 & {in3[6]});
 assign csa_tree_add_39_2_groupi_n_139 = (csa_tree_add_39_2_groupi_n_55 ^ {in3[6]});
 assign csa_tree_add_39_2_groupi_n_137 = (csa_tree_add_39_2_groupi_n_94 & csa_tree_add_39_2_groupi_n_59);
 assign csa_tree_add_39_2_groupi_n_140 = (csa_tree_add_39_2_groupi_n_94 ^ csa_tree_add_39_2_groupi_n_59);
 assign csa_tree_add_39_2_groupi_n_135 = ~(csa_tree_add_39_2_groupi_n_130 & ~csa_tree_add_39_2_groupi_n_120);
 assign csa_tree_add_39_2_groupi_n_134 = ~(csa_tree_add_39_2_groupi_n_10 & csa_tree_add_39_2_groupi_n_8);
 assign csa_tree_add_39_2_groupi_n_130 = ~(csa_tree_add_39_2_groupi_n_106 & csa_tree_add_39_2_groupi_n_20);
 assign csa_tree_add_39_2_groupi_n_129 = ~((csa_tree_add_39_2_groupi_n_30 & ~csa_tree_add_39_2_groupi_n_95)
    | ({in3[4]} & csa_tree_add_39_2_groupi_n_95));
 assign csa_tree_add_39_2_groupi_n_132 = (csa_tree_add_39_2_groupi_n_89 ^ {in3[3]});
 assign csa_tree_add_39_2_groupi_n_126 = ~(csa_tree_add_39_2_groupi_n_119 | ~csa_tree_add_39_2_groupi_n_105);
 assign csa_tree_add_39_2_groupi_n_125 = (csa_tree_add_39_2_groupi_n_97 ^ {in3[2]});
 assign csa_tree_add_39_2_groupi_n_122 = ~(({in3[7]} & ~csa_tree_add_39_2_groupi_n_99) | (csa_tree_add_39_2_groupi_n_38
    & csa_tree_add_39_2_groupi_n_99));
 assign csa_tree_add_39_2_groupi_n_121 = ~(({in3[1]} & ~csa_tree_add_39_2_groupi_n_66) | (csa_tree_add_39_2_groupi_n_29
    & csa_tree_add_39_2_groupi_n_66));
 assign csa_tree_add_39_2_groupi_n_120 = ~(csa_tree_add_39_2_groupi_n_58 | csa_tree_add_39_2_groupi_n_92);
 assign csa_tree_add_39_2_groupi_n_119 = ~(csa_tree_add_39_2_groupi_n_91 | ({in2[3]} & {in1[0]}));
 assign csa_tree_add_39_2_groupi_n_117 = ~(csa_tree_add_39_2_groupi_n_90 | csa_tree_add_39_2_groupi_n_93);
 assign csa_tree_add_39_2_groupi_n_112 = ~({in2[0]} & ({in1[3]} & {in3[3]}));
 assign csa_tree_add_39_2_groupi_n_111 = ~(csa_tree_add_39_2_groupi_n_66 | csa_tree_add_39_2_groupi_n_29);
 assign csa_tree_add_39_2_groupi_n_110 = ~(csa_tree_add_39_2_groupi_n_99 | csa_tree_add_39_2_groupi_n_38);
 assign csa_tree_add_39_2_groupi_n_107 = ~(csa_tree_add_39_2_groupi_n_63 & csa_tree_add_39_2_groupi_n_91);
 assign csa_tree_add_39_2_groupi_n_106 = ~(csa_tree_add_39_2_groupi_n_58 & csa_tree_add_39_2_groupi_n_92);
 assign csa_tree_add_39_2_groupi_n_105 = ~(csa_tree_add_39_2_groupi_n_91 & ~csa_tree_add_39_2_groupi_n_100);
 assign csa_tree_add_39_2_groupi_n_102 = ~(csa_tree_add_39_2_groupi_n_95 | csa_tree_add_39_2_groupi_n_30);
 assign csa_tree_add_39_2_groupi_n_101 = ~(csa_tree_add_39_2_groupi_n_96 | ~{in3[8]});
 assign csa_tree_add_39_2_groupi_n_89 = ~({in2[0]} & {in1[3]});
 assign csa_tree_add_39_2_groupi_n_88 = ({in2[4]} & {in1[7]});
 assign csa_tree_add_39_2_groupi_n_100 = ~({in2[3]} & {in1[0]});
 assign csa_tree_add_39_2_groupi_n_99 = ~({in2[0]} & {in1[7]});
 assign csa_tree_add_39_2_groupi_n_87 = ({in2[4]} & {in1[5]});
 assign csa_tree_add_39_2_groupi_n_98 = ~({in2[0]} & {in1[5]});
 assign csa_tree_add_39_2_groupi_n_97 = ~({in2[0]} & {in1[2]});
 assign csa_tree_add_39_2_groupi_n_86 = ({in2[3]} & {in1[7]});
 assign csa_tree_add_39_2_groupi_n_96 = ~({in2[1]} & {in1[7]});
 assign csa_tree_add_39_2_groupi_n_95 = ~({in2[0]} & {in1[4]});
 assign csa_tree_add_39_2_groupi_n_85 = ~(csa_tree_add_39_2_groupi_n_26 | csa_tree_add_39_2_groupi_n_27);
 assign csa_tree_add_39_2_groupi_n_94 = ~({in2[1]} & {in1[1]});
 assign csa_tree_add_39_2_groupi_n_93 = ~({in2[6]} & {in1[0]});
 assign csa_tree_add_39_2_groupi_n_84 = ~(csa_tree_add_39_2_groupi_n_34 | csa_tree_add_39_2_groupi_n_21);
 assign csa_tree_add_39_2_groupi_n_92 = ~({in2[2]} & {in1[2]});
 assign csa_tree_add_39_2_groupi_n_83 = ~(csa_tree_add_39_2_groupi_n_36 | csa_tree_add_39_2_groupi_n_37);
 assign csa_tree_add_39_2_groupi_n_82 = ({in2[5]} & {in1[6]});
 assign csa_tree_add_39_2_groupi_n_81 = ({in2[7]} & {in1[2]});
 assign csa_tree_add_39_2_groupi_n_80 = ~(csa_tree_add_39_2_groupi_n_24 | csa_tree_add_39_2_groupi_n_32);
 assign csa_tree_add_39_2_groupi_n_79 = ({in2[6]} & {in1[6]});
 assign csa_tree_add_39_2_groupi_n_78 = ~(csa_tree_add_39_2_groupi_n_25 | csa_tree_add_39_2_groupi_n_37);
 assign csa_tree_add_39_2_groupi_n_77 = ~(csa_tree_add_39_2_groupi_n_31 | csa_tree_add_39_2_groupi_n_32);
 assign csa_tree_add_39_2_groupi_n_76 = ~(csa_tree_add_39_2_groupi_n_26 | csa_tree_add_39_2_groupi_n_21);
 assign csa_tree_add_39_2_groupi_n_75 = ({in2[6]} & {in1[4]});
 assign csa_tree_add_39_2_groupi_n_91 = ~({in2[2]} & {in1[1]});
 assign csa_tree_add_39_2_groupi_n_90 = ~({in2[2]} & {in1[4]});
 assign csa_tree_add_39_2_groupi_n_74 = ~(csa_tree_add_39_2_groupi_n_36 | csa_tree_add_39_2_groupi_n_21);
 assign csa_tree_add_39_2_groupi_n_73 = ({in2[7]} & {in1[6]});
 assign csa_tree_add_39_2_groupi_n_72 = ({in2[7]} & {in1[5]});
 assign csa_tree_add_39_2_groupi_n_71 = ~(csa_tree_add_39_2_groupi_n_33 | csa_tree_add_39_2_groupi_n_22);
 assign csa_tree_add_39_2_groupi_n_70 = ~(csa_tree_add_39_2_groupi_n_34 | csa_tree_add_39_2_groupi_n_23);
 assign csa_tree_add_39_2_groupi_n_69 = ({in2[5]} & {in1[5]});
 assign csa_tree_add_39_2_groupi_n_65 = ~csa_tree_add_39_2_groupi_n_64;
 assign csa_tree_add_39_2_groupi_n_62 = ~csa_tree_add_39_2_groupi_n_63;
 assign csa_tree_add_39_2_groupi_n_68 = ~({in2[0]} & {in1[0]});
 assign csa_tree_add_39_2_groupi_n_57 = ~(csa_tree_add_39_2_groupi_n_36 | csa_tree_add_39_2_groupi_n_35);
 assign csa_tree_add_39_2_groupi_n_56 = ~(csa_tree_add_39_2_groupi_n_34 | csa_tree_add_39_2_groupi_n_35);
 assign csa_tree_add_39_2_groupi_n_55 = ~(csa_tree_add_39_2_groupi_n_25 | csa_tree_add_39_2_groupi_n_22);
 assign csa_tree_add_39_2_groupi_n_54 = ~(csa_tree_add_39_2_groupi_n_34 | csa_tree_add_39_2_groupi_n_37);
 assign csa_tree_add_39_2_groupi_n_67 = ~(csa_tree_add_39_2_groupi_n_33 | csa_tree_add_39_2_groupi_n_27);
 assign csa_tree_add_39_2_groupi_n_66 = ~({in2[1]} & {in1[0]});
 assign csa_tree_add_39_2_groupi_n_53 = ~(csa_tree_add_39_2_groupi_n_26 | csa_tree_add_39_2_groupi_n_23);
 assign csa_tree_add_39_2_groupi_n_52 = ~(csa_tree_add_39_2_groupi_n_31 | csa_tree_add_39_2_groupi_n_22);
 assign csa_tree_add_39_2_groupi_n_51 = ~(csa_tree_add_39_2_groupi_n_26 | csa_tree_add_39_2_groupi_n_22);
 assign csa_tree_add_39_2_groupi_n_64 = ~({in2[3]} & {in1[3]});
 assign csa_tree_add_39_2_groupi_n_50 = ~(csa_tree_add_39_2_groupi_n_36 | csa_tree_add_39_2_groupi_n_23);
 assign csa_tree_add_39_2_groupi_n_63 = ~({in2[1]} & {in1[2]});
 assign csa_tree_add_39_2_groupi_n_49 = ~(csa_tree_add_39_2_groupi_n_36 | csa_tree_add_39_2_groupi_n_32);
 assign csa_tree_add_39_2_groupi_n_48 = ~(csa_tree_add_39_2_groupi_n_34 | csa_tree_add_39_2_groupi_n_27);
 assign csa_tree_add_39_2_groupi_n_47 = ~(csa_tree_add_39_2_groupi_n_33 | csa_tree_add_39_2_groupi_n_32);
 assign csa_tree_add_39_2_groupi_n_61 = ~(csa_tree_add_39_2_groupi_n_31 | csa_tree_add_39_2_groupi_n_23);
 assign csa_tree_add_39_2_groupi_n_46 = ~(csa_tree_add_39_2_groupi_n_28 | csa_tree_add_39_2_groupi_n_27);
 assign csa_tree_add_39_2_groupi_n_45 = ({in2[7]} & {in1[7]});
 assign csa_tree_add_39_2_groupi_n_44 = ~(csa_tree_add_39_2_groupi_n_24 | csa_tree_add_39_2_groupi_n_22);
 assign csa_tree_add_39_2_groupi_n_60 = ~({in2[3]} & {in1[2]});
 assign csa_tree_add_39_2_groupi_n_59 = ~({in2[2]} & {in1[0]});
 assign csa_tree_add_39_2_groupi_n_43 = ~(csa_tree_add_39_2_groupi_n_24 | csa_tree_add_39_2_groupi_n_27);
 assign csa_tree_add_39_2_groupi_n_42 = ~({in2[4]} & {in1[0]});
 assign csa_tree_add_39_2_groupi_n_58 = ~({in2[1]} & {in1[3]});
 assign csa_tree_add_39_2_groupi_n_41 = ~(csa_tree_add_39_2_groupi_n_31 | csa_tree_add_39_2_groupi_n_35);
 assign csa_tree_add_39_2_groupi_n_40 = ~(csa_tree_add_39_2_groupi_n_28 | csa_tree_add_39_2_groupi_n_23);
 assign csa_tree_add_39_2_groupi_n_39 = ~(csa_tree_add_39_2_groupi_n_28 | csa_tree_add_39_2_groupi_n_37);
 assign csa_tree_add_39_2_groupi_n_38 = ~{in3[7]};
 assign csa_tree_add_39_2_groupi_n_37 = ~{in1[1]};
 assign csa_tree_add_39_2_groupi_n_36 = ~{in2[6]};
 assign csa_tree_add_39_2_groupi_n_35 = ~{in1[7]};
 assign csa_tree_add_39_2_groupi_n_34 = ~{in2[5]};
 assign csa_tree_add_39_2_groupi_n_33 = ~{in2[1]};
 assign csa_tree_add_39_2_groupi_n_32 = ~{in1[5]};
 assign csa_tree_add_39_2_groupi_n_31 = ~{in2[2]};
 assign csa_tree_add_39_2_groupi_n_30 = ~{in3[4]};
 assign csa_tree_add_39_2_groupi_n_29 = ~{in3[1]};
 assign csa_tree_add_39_2_groupi_n_28 = ~{in2[7]};
 assign csa_tree_add_39_2_groupi_n_27 = ~{in1[4]};
 assign csa_tree_add_39_2_groupi_n_26 = ~{in2[4]};
 assign csa_tree_add_39_2_groupi_n_25 = ~{in2[0]};
 assign csa_tree_add_39_2_groupi_n_24 = ~{in2[3]};
 assign csa_tree_add_39_2_groupi_n_23 = ~{in1[3]};
 assign csa_tree_add_39_2_groupi_n_22 = ~{in1[6]};
 assign csa_tree_add_39_2_groupi_n_21 = ~{in1[2]};
 assign csa_tree_add_39_2_groupi_n_19 = ({in2[5]} & {in1[0]});
 assign csa_tree_add_39_2_groupi_n_18 = ({in2[4]} & {in1[1]});
 assign csa_tree_add_39_2_groupi_n_17 = ~(csa_tree_add_39_2_groupi_n_208 & ~n_106);
 assign csa_tree_add_39_2_groupi_n_16 = (csa_tree_add_39_2_groupi_n_191 ^ csa_tree_add_39_2_groupi_n_184);
 assign csa_tree_add_39_2_groupi_n_15 = ~(n_109 & ~csa_tree_add_39_2_groupi_n_182);
 assign csa_tree_add_39_2_groupi_n_14 = ~(csa_tree_add_39_2_groupi_n_4 ^ csa_tree_add_39_2_groupi_n_134);
 assign csa_tree_add_39_2_groupi_n_12 = ~(csa_tree_add_39_2_groupi_n_132 ^ csa_tree_add_39_2_groupi_n_1);
 assign csa_tree_add_39_2_groupi_n_10 = ~(csa_tree_add_39_2_groupi_n_107 & ~csa_tree_add_39_2_groupi_n_100);
 assign csa_tree_add_39_2_groupi_n_9 = (csa_tree_add_39_2_groupi_n_94 | csa_tree_add_39_2_groupi_n_59);
 assign csa_tree_add_39_2_groupi_n_8 = ~(csa_tree_add_39_2_groupi_n_62 & ~csa_tree_add_39_2_groupi_n_91);
 assign csa_tree_add_39_2_groupi_n_7 = (n_114 ^ csa_tree_add_39_2_groupi_n_67);
 assign csa_tree_add_39_2_groupi_n_6 = ~(csa_tree_add_39_2_groupi_n_60 & ~csa_tree_add_39_2_groupi_n_61);
 assign csa_tree_add_39_2_groupi_n_5 = ~(csa_tree_add_39_2_groupi_n_61 & ~csa_tree_add_39_2_groupi_n_60);
 assign csa_tree_add_39_2_groupi_n_4 = ~(n_116 ^ csa_tree_add_39_2_groupi_n_58);
 assign csa_tree_add_39_2_groupi_n_3 = ~(csa_tree_add_39_2_groupi_n_68 | ~{in3[0]});
 assign csa_tree_add_39_2_groupi_n_2 = ~(csa_tree_add_39_2_groupi_n_28 | ~{in1[0]});
 assign csa_tree_add_39_2_groupi_n_1 = ~(csa_tree_add_39_2_groupi_n_97 | ~{in3[2]});
 assign csa_tree_add_39_2_groupi_n_0 = ~(csa_tree_add_39_2_groupi_n_98 | ~{in3[5]});
 assign n_54 = ~csa_tree_add_39_2_groupi_n_301;
 assign csa_tree_add_39_2_groupi_n_301 = ((csa_tree_add_39_2_groupi_n_195 & n_57) | ((n_57 & {in3[15]})
    | ({in3[15]} & csa_tree_add_39_2_groupi_n_195)));
 assign n_55 = (n_57 ^ ({in3[15]} ^ csa_tree_add_39_2_groupi_n_195));
 assign n_57 = ((csa_tree_add_39_2_groupi_n_251 & n_59) | ((n_59 & csa_tree_add_39_2_groupi_n_196) |
    (csa_tree_add_39_2_groupi_n_196 & csa_tree_add_39_2_groupi_n_251)));
 assign n_56 = (n_59 ^ (csa_tree_add_39_2_groupi_n_196 ^ csa_tree_add_39_2_groupi_n_251));
 assign n_59 = ((csa_tree_add_39_2_groupi_n_266 & n_61) | ((n_61 & csa_tree_add_39_2_groupi_n_252) |
    (csa_tree_add_39_2_groupi_n_252 & csa_tree_add_39_2_groupi_n_266)));
 assign n_58 = (n_61 ^ (csa_tree_add_39_2_groupi_n_252 ^ csa_tree_add_39_2_groupi_n_266));
 assign n_61 = ((csa_tree_add_39_2_groupi_n_268 & n_63) | ((n_63 & csa_tree_add_39_2_groupi_n_267) |
    (csa_tree_add_39_2_groupi_n_267 & csa_tree_add_39_2_groupi_n_268)));
 assign n_60 = (n_63 ^ (csa_tree_add_39_2_groupi_n_267 ^ csa_tree_add_39_2_groupi_n_268));
 assign n_63 = ((csa_tree_add_39_2_groupi_n_269 & n_65) | ((n_65 & csa_tree_add_39_2_groupi_n_278) |
    (csa_tree_add_39_2_groupi_n_278 & csa_tree_add_39_2_groupi_n_269)));
 assign n_62 = (n_65 ^ (csa_tree_add_39_2_groupi_n_278 ^ csa_tree_add_39_2_groupi_n_269));
 assign n_65 = ((csa_tree_add_39_2_groupi_n_279 & n_67) | ((n_67 & csa_tree_add_39_2_groupi_n_280) |
    (csa_tree_add_39_2_groupi_n_280 & csa_tree_add_39_2_groupi_n_279)));
 assign n_64 = (n_67 ^ (csa_tree_add_39_2_groupi_n_280 ^ csa_tree_add_39_2_groupi_n_279));
 assign n_67 = ((csa_tree_add_39_2_groupi_n_281 & n_69) | ((n_69 & csa_tree_add_39_2_groupi_n_274) |
    (csa_tree_add_39_2_groupi_n_274 & csa_tree_add_39_2_groupi_n_281)));
 assign n_66 = (n_69 ^ (csa_tree_add_39_2_groupi_n_274 ^ csa_tree_add_39_2_groupi_n_281));
 assign n_69 = ((csa_tree_add_39_2_groupi_n_275 & n_71) | ((n_71 & csa_tree_add_39_2_groupi_n_272) |
    (csa_tree_add_39_2_groupi_n_272 & csa_tree_add_39_2_groupi_n_275)));
 assign n_68 = (n_71 ^ (csa_tree_add_39_2_groupi_n_272 ^ csa_tree_add_39_2_groupi_n_275));
 assign n_71 = ((n_73 & csa_tree_add_39_2_groupi_n_273) | ((csa_tree_add_39_2_groupi_n_273 & csa_tree_add_39_2_groupi_n_265)
    | (csa_tree_add_39_2_groupi_n_265 & n_73)));
 assign n_70 = (csa_tree_add_39_2_groupi_n_273 ^ (csa_tree_add_39_2_groupi_n_265 ^ n_73));
 assign n_73 = ((n_75 & n_102) | ((n_102 & csa_tree_add_39_2_groupi_n_247) | (csa_tree_add_39_2_groupi_n_247
    & n_75)));
 assign n_72 = (n_102 ^ (csa_tree_add_39_2_groupi_n_247 ^ n_75));
 assign n_75 = ((n_104 & n_77) | ((n_77 & csa_tree_add_39_2_groupi_n_221) | (csa_tree_add_39_2_groupi_n_221
    & n_104)));
 assign n_74 = (n_77 ^ (csa_tree_add_39_2_groupi_n_221 ^ n_104));
 assign {out1[31]} = ~(n_80 ^ n_48);
 assign n_77 = ((n_79 & n_107) | ((n_107 & csa_tree_add_39_2_groupi_n_190) | (csa_tree_add_39_2_groupi_n_190
    & n_79)));
 assign n_76 = (n_107 ^ (csa_tree_add_39_2_groupi_n_190 ^ n_79));
 assign {out1[30]} = ~(n_81 ^ n_47);
 assign n_80 = ~(n_47 & ~n_81);
 assign n_79 = ((n_84 & n_108) | ((n_108 & csa_tree_add_39_2_groupi_n_154) | (csa_tree_add_39_2_groupi_n_154
    & n_84)));
 assign n_78 = (n_108 ^ (csa_tree_add_39_2_groupi_n_154 ^ n_84));
 assign {out1[29]} = ~(n_82 ^ n_50);
 assign n_81 = ~(n_50 & ~n_82);
 assign {out1[28]} = ~(n_85 ^ n_49);
 assign n_82 = ~(n_49 & ~n_85);
 assign n_84 = ((n_2 & n_110) | ((n_110 & csa_tree_add_39_2_groupi_n_111) | (csa_tree_add_39_2_groupi_n_111
    & n_2)));
 assign n_83 = (n_110 ^ (csa_tree_add_39_2_groupi_n_111 ^ n_2));
 assign {out1[27]} = ~(n_0 ^ n_51);
 assign n_85 = ~(n_51 & ~n_0);
 assign {out1[26]} = ~(n_53 ^ n_52);
 assign n_2 = ((csa_tree_add_39_2_groupi_n_78 & csa_tree_add_39_2_groupi_n_121) | ((csa_tree_add_39_2_groupi_n_121
    & csa_tree_add_39_2_groupi_n_3) | (csa_tree_add_39_2_groupi_n_3 & csa_tree_add_39_2_groupi_n_78)));
 assign n_1 = (csa_tree_add_39_2_groupi_n_121 ^ (csa_tree_add_39_2_groupi_n_3 ^ csa_tree_add_39_2_groupi_n_78));
 assign n_0 = ~(n_52 & ~n_53);
 assign n_9 = ~(csa_tree_add_39_2_groupi_n_316 ^ {in3[24]});
 assign n_8 = ~(csa_tree_add_39_2_groupi_n_318 ^ {in3[25]});
 assign n_11 = ~(csa_tree_add_39_2_groupi_n_68 ^ {in3[0]});
 assign n_12 = ~(csa_tree_add_39_2_groupi_n_314 ^ {in3[23]});
 assign n_5 = ~(csa_tree_add_39_2_groupi_n_312 ^ {in3[22]});
 assign n_4 = ~(csa_tree_add_39_2_groupi_n_306 ^ {in3[19]});
 assign n_3 = ~(csa_tree_add_39_2_groupi_n_308 ^ {in3[20]});
 assign n_6 = ~(csa_tree_add_39_2_groupi_n_310 ^ {in3[21]});
 assign n_7 = ~(csa_tree_add_39_2_groupi_n_304 ^ {in3[18]});
 assign n_10 = ~(csa_tree_add_39_2_groupi_n_302 ^ {in3[17]});
 assign n_13 = ~({in3[25]} & ~csa_tree_add_39_2_groupi_n_318);
 assign n_102 = ~(n_103 ^ csa_tree_add_39_2_groupi_n_16);
 assign n_103 = ~(csa_tree_add_39_2_groupi_n_218 ^ csa_tree_add_39_2_groupi_n_222);
 assign n_104 = ~(n_106 ^ n_105);
 assign n_105 = ~(csa_tree_add_39_2_groupi_n_185 ^ csa_tree_add_39_2_groupi_n_201);
 assign n_106 = (csa_tree_add_39_2_groupi_n_199 ^ csa_tree_add_39_2_groupi_n_7);
 assign n_107 = ~(csa_tree_add_39_2_groupi_n_14 ^ csa_tree_add_39_2_groupi_n_202);
 assign n_108 = ~(n_111 ^ csa_tree_add_39_2_groupi_n_12);
 assign n_109 = ((csa_tree_add_39_2_groupi_n_65 & ~n_115) | (csa_tree_add_39_2_groupi_n_64 & n_115));
 assign n_110 = ~(csa_tree_add_39_2_groupi_n_140 ^ csa_tree_add_39_2_groupi_n_125);
 assign n_111 = ((csa_tree_add_39_2_groupi_n_62 & ~csa_tree_add_39_2_groupi_n_126) | (csa_tree_add_39_2_groupi_n_63
    & csa_tree_add_39_2_groupi_n_126));
 assign n_112 = ~(csa_tree_add_39_2_groupi_n_96 ^ {in3[8]});
 assign n_113 = ~(csa_tree_add_39_2_groupi_n_98 ^ {in3[5]});
 assign n_114 = (csa_tree_add_39_2_groupi_n_61 ^ csa_tree_add_39_2_groupi_n_60);
 assign n_115 = ~(csa_tree_add_39_2_groupi_n_90 ^ csa_tree_add_39_2_groupi_n_93);
 assign n_116 = (csa_tree_add_39_2_groupi_n_20 ^ csa_tree_add_39_2_groupi_n_92);
endmodule
