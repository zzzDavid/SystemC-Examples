`timescale 1ps / 1ps
module dut_Div_64Ux2U_32U_4(
          in2,
          in1,
          out1,
          clk,
          stall
);
   input [63:0] in2;
   input [1:0] in1;
   output [31:0] out1;
   input clk;
   input stall;
wire sub_289_2_n_1, sub_289_2_n_2, sub_308_2_n_0, sub_308_2_n_1, sub_308_2_n_2,
     sub_308_2_n_3, sub_308_2_n_4, sub_308_2_n_6, sub_327_2_n_1, sub_327_2_n_2,
     sub_327_2_n_3, sub_327_2_n_4, sub_327_2_n_5, sub_327_2_n_7, sub_327_2_n_9,
     sub_346_2_n_1, sub_346_2_n_2, sub_346_2_n_3, sub_346_2_n_4, sub_346_2_n_6,
     sub_346_2_n_7, sub_346_2_n_9, sub_365_2_n_0, sub_365_2_n_2, sub_365_2_n_3,
     sub_365_2_n_5, sub_384_2_n_0, sub_384_2_n_1, sub_384_2_n_2, sub_384_2_n_4,
     sub_403_2_n_0, sub_403_2_n_1, sub_403_2_n_2, sub_403_2_n_4, sub_422_2_n_0,
     sub_422_2_n_2, sub_422_2_n_3, sub_422_2_n_5, sub_441_2_n_0, sub_441_2_n_1,
     sub_441_2_n_2, sub_441_2_n_4, sub_460_2_n_0, sub_460_2_n_1, sub_460_2_n_2,
     sub_460_2_n_4, sub_479_2_n_0, sub_479_2_n_1, sub_479_2_n_2, sub_479_2_n_5,
     sub_479_2_n_6, sub_498_2_n_0, sub_498_2_n_1, sub_498_2_n_2, sub_498_2_n_4,
     sub_517_2_n_0, sub_517_2_n_1, sub_517_2_n_2, sub_517_2_n_4, sub_536_2_n_0,
     sub_536_2_n_2, sub_536_2_n_3, sub_536_2_n_5, sub_555_2_n_0, sub_555_2_n_1,
     sub_555_2_n_2, sub_555_2_n_4, sub_574_2_n_0, sub_574_2_n_1, sub_574_2_n_2,
     sub_574_2_n_4, sub_593_2_n_0, sub_593_2_n_2, sub_593_2_n_3, sub_593_2_n_5,
     sub_612_2_n_0, sub_612_2_n_1, sub_612_2_n_2, sub_612_2_n_4, sub_631_2_n_0,
     sub_631_2_n_2, sub_631_2_n_3, sub_631_2_n_5, sub_650_2_n_0, sub_650_2_n_1,
     sub_650_2_n_2, sub_650_2_n_4, sub_669_2_n_0, sub_669_2_n_2, sub_669_2_n_3,
     sub_669_2_n_5, sub_688_2_n_0, sub_688_2_n_1, sub_688_2_n_2, sub_688_2_n_3,
     sub_688_2_n_5, sub_688_2_n_6, sub_688_2_n_8, sub_707_2_n_0, sub_707_2_n_2,
     sub_707_2_n_3, sub_707_2_n_5, sub_726_2_n_0, sub_726_2_n_1, sub_726_2_n_2,
     sub_726_2_n_3, sub_726_2_n_5, sub_726_2_n_6, sub_726_2_n_8, sub_745_2_n_0,
     sub_745_2_n_2, sub_745_2_n_3, sub_745_2_n_5, sub_764_2_n_0, sub_764_2_n_1,
     sub_764_2_n_2, sub_764_2_n_3, sub_764_2_n_5, sub_764_2_n_6, sub_764_2_n_8,
     sub_783_2_n_0, sub_783_2_n_2, sub_783_2_n_3, sub_783_2_n_5, sub_802_2_n_1,
     sub_802_2_n_2, sub_802_2_n_3, sub_802_2_n_4, sub_802_2_n_6, sub_802_2_n_7,
     sub_802_2_n_9, sub_821_2_n_1, sub_821_2_n_2, sub_821_2_n_3, sub_821_2_n_4,
     sub_821_2_n_6, sub_821_2_n_7, sub_821_2_n_9, sub_840_2_n_1, sub_840_2_n_2,
     sub_840_2_n_3, sub_840_2_n_4, sub_840_2_n_6, sub_840_2_n_7, sub_840_2_n_9,
     sub_859_2_n_1, sub_859_2_n_2, sub_859_2_n_3, sub_859_2_n_4, sub_859_2_n_6,
     sub_859_2_n_7, sub_859_2_n_9, sub_878_2_n_1, sub_878_2_n_2, sub_878_2_n_3,
     sub_878_2_n_4, sub_878_2_n_6, sub_878_2_n_7, sub_878_2_n_9, sub_897_2_n_1,
     sub_897_2_n_2, sub_897_2_n_3, sub_897_2_n_4, sub_897_2_n_6, sub_897_2_n_7,
     sub_897_2_n_9, sub_918_2_n_1, sub_918_2_n_2, sub_918_2_n_3, sub_918_2_n_4,
     sub_918_2_n_6, sub_918_2_n_7, sub_918_2_n_9, sub_939_2_n_1, sub_939_2_n_2,
     sub_939_2_n_3, sub_939_2_n_4, sub_939_2_n_6, sub_939_2_n_7, sub_939_2_n_9,
     sub_960_2_n_1, sub_960_2_n_2, sub_960_2_n_3, sub_960_2_n_4, sub_960_2_n_6,
     sub_960_2_n_7, sub_960_2_n_9, sub_981_2_n_1, sub_981_2_n_2, sub_981_2_n_3,
     sub_981_2_n_4, sub_981_2_n_6, sub_981_2_n_7, sub_981_2_n_9, sub_1002_2_n_1,
     sub_1002_2_n_2, sub_1002_2_n_3, sub_1002_2_n_4, sub_1002_2_n_6,
     sub_1002_2_n_7, sub_1002_2_n_9, sub_1023_2_n_1, sub_1023_2_n_2,
     sub_1023_2_n_3, sub_1023_2_n_4, sub_1023_2_n_6, sub_1023_2_n_7,
     sub_1023_2_n_9, sub_1044_2_n_1, sub_1044_2_n_2, sub_1044_2_n_3,
     sub_1044_2_n_4, sub_1044_2_n_6, sub_1044_2_n_7, sub_1044_2_n_9,
     sub_1065_2_n_1, sub_1065_2_n_2, sub_1065_2_n_3, sub_1065_2_n_4,
     sub_1065_2_n_6, sub_1065_2_n_7, sub_1065_2_n_9, sub_1086_2_n_1,
     sub_1086_2_n_2, sub_1086_2_n_3, sub_1086_2_n_4, sub_1086_2_n_6,
     sub_1086_2_n_7, sub_1086_2_n_9, sub_1107_2_n_1, sub_1107_2_n_2,
     sub_1107_2_n_3, sub_1107_2_n_4, sub_1107_2_n_6, sub_1107_2_n_7,
     sub_1107_2_n_9, sub_1128_2_n_2, sub_1128_2_n_5, sub_1149_2_n_1,
     sub_1149_2_n_2, sub_1149_2_n_4, sub_1170_2_n_2, sub_1170_2_n_4,
     sub_1191_2_n_2, sub_1191_2_n_4, sub_1212_2_n_1, sub_1212_2_n_2,
     sub_1212_2_n_4, sub_1233_2_n_1, sub_1233_2_n_2, sub_1233_2_n_4,
     sub_1254_2_n_1, sub_1254_2_n_2, sub_1254_2_n_4, sub_1275_2_n_1,
     sub_1275_2_n_2, sub_1275_2_n_4, sub_1296_2_n_1, sub_1296_2_n_2,
     sub_1296_2_n_4, sub_1317_2_n_1, sub_1317_2_n_2, sub_1317_2_n_4,
     sub_1338_2_n_1, sub_1338_2_n_2, sub_1338_2_n_4, sub_1359_2_n_1,
     sub_1359_2_n_2, sub_1359_2_n_4, sub_1380_2_n_1, sub_1380_2_n_2,
     sub_1380_2_n_4, sub_1401_2_n_1, sub_1401_2_n_2, sub_1401_2_n_4,
     sub_1422_2_n_1, sub_1422_2_n_2, sub_1422_2_n_4, sub_1443_2_n_1,
     sub_1443_2_n_2, sub_1443_2_n_4, sub_1464_2_n_1, sub_1464_2_n_2,
     sub_1464_2_n_4, sub_1485_2_n_1, sub_1485_2_n_2, sub_1485_2_n_4,
     sub_1506_2_n_1, sub_1506_2_n_2, sub_1506_2_n_4, sub_1527_2_n_1,
     sub_1527_2_n_2, sub_1527_2_n_4, sub_1546_2_n_1, sub_1546_2_n_4, n_0, n_1,
     n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15,
     n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_27,
     n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39,
     n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51,
     n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63,
     n_64, n_65, n_67, n_68, clk, stall, n_106, n_107, n_108, n_109, n_110,
     n_111, n_112, n_115, n_116, n_117, n_120, n_121, n_122, n_123, n_125, n_126,
     n_127, n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137,
     n_138, n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149,
     n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160,
     n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_170, n_171, n_172,
     n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183,
     n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193, n_195, n_196,
     n_197, n_198, n_199, n_200, n_201, n_202, n_205, n_206, n_207, n_208, n_209,
     n_210, n_211, n_212, n_215, n_216, n_217, n_218, n_219, n_220, n_221, n_222,
     n_225, n_226, n_227, n_229, n_230, n_231, n_232, n_235, n_236, n_237, n_240,
     n_241, n_242, n_245, n_246, n_247, n_250, n_251, n_252, n_255, n_256, n_257,
     n_260, n_261, n_262, n_265, n_266, n_267, n_268, n_269, n_270, n_271, n_274,
     n_275, n_276, n_279, n_280, n_281, n_283, n_284, n_285, n_286, n_288, n_289,
     n_290, n_291, n_293, n_294, n_295, n_296, n_298, n_299, n_300, n_303, n_304,
     n_305, n_308, n_309, n_310, n_311, n_313, n_314, n_315, n_319, n_320, n_321,
     n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330, n_331, n_332,
     n_333, n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341, n_342, n_343,
     n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352, n_353, n_354,
     n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363, n_364, n_365,
     n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376,
     n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385, n_386, n_387,
     n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395, n_396, n_397, n_398,
     n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_430, n_431, n_432, n_433,
     n_434, n_437, n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446,
     n_447, n_448, n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457,
     n_458, n_459, n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468,
     n_469, n_470, n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479,
     n_480, n_481, n_482, n_483, in2_190_2_;
 reg out1_0_L0_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         out1_0_L0_reg_N30 <= n_479;
 assign n_0 = out1_0_L0_reg_N30;
 reg retime_s1_1_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_1_reg_reg_N30 <= {in1[0]};
 assign n_1 = retime_s1_1_reg_reg_N30;
 reg retime_s1_2_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_2_reg_reg_N30 <= {in2[1]};
 assign n_2 = retime_s1_2_reg_reg_N30;
 reg retime_s1_3_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_3_reg_reg_N30 <= n_65;
 assign n_267 = retime_s1_3_reg_reg_N30;
 reg retime_s1_4_reg_reg_N30;
 always @(posedge clk)
         retime_s1_4_reg_reg_N30 <= n_34;
 assign sub_1149_2_n_1 = retime_s1_4_reg_reg_N30;
 reg retime_s1_5_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_5_reg_reg_N30 <= {in2[11]};
 assign n_3 = retime_s1_5_reg_reg_N30;
 reg retime_s1_6_reg_reg_N30;
 always @(posedge clk)
         retime_s1_6_reg_reg_N30 <= n_47;
 assign n_4 = retime_s1_6_reg_reg_N30;
 reg retime_s1_7_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_7_reg_reg_N30 <= {in2[17]};
 assign n_5 = retime_s1_7_reg_reg_N30;
 reg retime_s1_8_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_8_reg_reg_N30 <= {in2[3]};
 assign n_6 = retime_s1_8_reg_reg_N30;
 reg retime_s1_9_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_9_reg_reg_N30 <= {in2[23]};
 assign n_7 = retime_s1_9_reg_reg_N30;
 reg retime_s1_10_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_10_reg_reg_N30 <= {in2[15]};
 assign n_8 = retime_s1_10_reg_reg_N30;
 reg retime_s1_11_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_11_reg_reg_N30 <= {in2[29]};
 assign n_9 = retime_s1_11_reg_reg_N30;
 reg retime_s1_12_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_12_reg_reg_N30 <= {in2[18]};
 assign n_10 = retime_s1_12_reg_reg_N30;
 reg retime_s1_13_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_13_reg_reg_N30 <= {in2[9]};
 assign n_11 = retime_s1_13_reg_reg_N30;
 reg retime_s1_14_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_14_reg_reg_N30 <= {in2[20]};
 assign n_12 = retime_s1_14_reg_reg_N30;
 reg retime_s1_15_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_15_reg_reg_N30 <= {in2[4]};
 assign n_13 = retime_s1_15_reg_reg_N30;
 reg retime_s1_16_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_16_reg_reg_N30 <= {in2[10]};
 assign n_14 = retime_s1_16_reg_reg_N30;
 reg retime_s1_17_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_17_reg_reg_N30 <= {in2[21]};
 assign n_15 = retime_s1_17_reg_reg_N30;
 reg retime_s1_18_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_18_reg_reg_N30 <= {in2[25]};
 assign n_16 = retime_s1_18_reg_reg_N30;
 reg retime_s1_19_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_19_reg_reg_N30 <= {in2[22]};
 assign n_17 = retime_s1_19_reg_reg_N30;
 reg retime_s1_20_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_20_reg_reg_N30 <= {in2[26]};
 assign n_18 = retime_s1_20_reg_reg_N30;
 reg retime_s1_21_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_21_reg_reg_N30 <= {in2[24]};
 assign n_19 = retime_s1_21_reg_reg_N30;
 reg retime_s1_22_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_22_reg_reg_N30 <= {in2[19]};
 assign n_20 = retime_s1_22_reg_reg_N30;
 reg retime_s1_23_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_23_reg_reg_N30 <= {in2[2]};
 assign n_21 = retime_s1_23_reg_reg_N30;
 reg retime_s1_24_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_24_reg_reg_N30 <= {in2[16]};
 assign n_22 = retime_s1_24_reg_reg_N30;
 reg retime_s1_25_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_25_reg_reg_N30 <= {in2[14]};
 assign n_23 = retime_s1_25_reg_reg_N30;
 reg retime_s1_26_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_26_reg_reg_N30 <= {in2[7]};
 assign n_24 = retime_s1_26_reg_reg_N30;
 reg retime_s1_27_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_27_reg_reg_N30 <= {in2[8]};
 assign n_25 = retime_s1_27_reg_reg_N30;
 reg retime_s1_28_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_28_reg_reg_N30 <= {in2[13]};
 assign n_26 = retime_s1_28_reg_reg_N30;
 reg retime_s1_29_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_29_reg_reg_N30 <= {in2[12]};
 assign n_27 = retime_s1_29_reg_reg_N30;
 reg retime_s1_30_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_30_reg_reg_N30 <= {in2[5]};
 assign n_28 = retime_s1_30_reg_reg_N30;
 reg retime_s1_31_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_31_reg_reg_N30 <= {in2[27]};
 assign n_29 = retime_s1_31_reg_reg_N30;
 reg retime_s1_32_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_32_reg_reg_N30 <= n_454;
 assign n_30 = retime_s1_32_reg_reg_N30;
 reg retime_s1_33_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_33_reg_reg_N30 <= {in2[28]};
 assign n_31 = retime_s1_33_reg_reg_N30;
 reg retime_s1_34_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_34_reg_reg_N30 <= {in2[6]};
 assign n_32 = retime_s1_34_reg_reg_N30;
 reg retime_s1_35_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_35_reg_reg_N30 <= {in2[30]};
 assign n_33 = retime_s1_35_reg_reg_N30;
 assign n_218 = ((n_216 & ~n_471) | ({in2[41]} & n_471));
 assign n_208 = ((n_206 & ~n_470) | ({in2[43]} & n_470));
 assign n_198 = ((n_196 & ~n_469) | ({in2[45]} & n_469));
 assign n_193 = ((n_191 & ~n_189) | ({in2[46]} & n_189));
 assign n_188 = ((n_186 & ~n_468) | ({in2[47]} & n_468));
 assign n_183 = ((n_181 & ~n_179) | ({in2[48]} & n_179));
 assign n_178 = ((n_176 & ~n_174) | ({in2[49]} & n_174));
 assign n_173 = ((n_171 & ~n_467) | ({in2[50]} & n_467));
 assign n_168 = ((n_166 & ~n_164) | ({in2[51]} & n_164));
 assign n_163 = ((n_161 & ~n_159) | ({in2[52]} & n_159));
 assign n_158 = ((n_156 & ~n_154) | ({in2[53]} & n_154));
 assign n_153 = ((n_151 & ~n_149) | ({in2[54]} & n_149));
 assign n_148 = ((n_146 & ~n_144) | ({in2[55]} & n_144));
 assign n_143 = ((n_141 & ~n_466) | ({in2[56]} & n_466));
 assign n_138 = ((n_136 & ~n_134) | ({in2[57]} & n_134));
 assign n_108 = ~(n_431 & n_430);
 assign n_430 = ~(n_106 & {in2[63]});
 assign n_431 = ~(n_432 & n_107);
 assign n_432 = ~n_106;
 assign n_123 = ~((n_434 & ~n_464) | (n_433 & n_464));
 assign n_433 = ~{in2[60]};
 assign n_434 = ~n_121;
 assign {out1[20]} = ~n_483;
 assign {out1[21]} = ~n_313;
 assign {out1[22]} = ~n_308;
 assign {out1[23]} = ~n_303;
 assign {out1[24]} = ~n_298;
 assign {out1[25]} = ~n_293;
 assign {out1[26]} = ~n_288;
 assign {out1[27]} = ~n_283;
 assign {out1[28]} = ~n_481;
 assign {out1[29]} = ~n_480;
 assign {out1[15]} = ~n_338;
 assign {out1[0]} = ~in2_190_2_;
 assign n_262 = ((n_260 & ~n_478) | (n_440 & n_478));
 assign n_276 = ((n_274 & ~n_480) | (n_452 & n_480));
 assign n_257 = ((n_255 & ~n_477) | (n_441 & n_477));
 assign n_281 = ((n_279 & ~n_481) | (n_459 & n_481));
 assign n_252 = ((n_250 & ~n_476) | (n_442 & n_476));
 assign n_286 = ((n_284 & ~n_283) | (n_457 & n_283));
 assign n_247 = ((n_245 & ~n_475) | (n_443 & n_475));
 assign n_291 = ((n_289 & ~n_288) | (n_456 & n_288));
 assign n_242 = ((n_240 & ~n_474) | (n_444 & n_474));
 assign n_296 = ((n_294 & ~n_293) | (n_455 & n_293));
 assign n_237 = ((n_235 & ~n_473) | (n_446 & n_473));
 assign n_232 = ((n_230 & ~n_229) | (n_448 & n_229));
 assign n_227 = ((n_225 & ~n_472) | (n_449 & n_472));
 assign n_311 = ((n_309 & ~n_308) | (n_458 & n_308));
 assign n_222 = ((n_220 & ~n_219) | (n_218 & n_219));
 assign n_217 = ((n_215 & ~n_471) | (n_437 & n_471));
 assign n_320 = ((n_319 & ~n_483) | (n_453 & n_483));
 assign n_212 = ((n_210 & ~n_209) | (n_208 & n_209));
 assign n_324 = ((n_323 & ~n_322) | (n_321 & n_322));
 assign n_207 = ((n_205 & ~n_470) | (n_438 & n_470));
 assign n_328 = ((n_327 & ~n_326) | (n_325 & n_326));
 assign n_202 = ((n_200 & ~n_199) | (n_198 & n_199));
 assign n_332 = ((n_331 & ~n_330) | (n_329 & n_330));
 assign n_197 = ((n_195 & ~n_469) | (n_193 & n_469));
 assign n_336 = ((n_335 & ~n_334) | (n_333 & n_334));
 assign n_192 = ((n_190 & ~n_189) | (n_188 & n_189));
 assign n_340 = ((n_339 & ~n_338) | (n_337 & n_338));
 assign n_187 = ((n_185 & ~n_468) | (n_183 & n_468));
 assign n_345 = ((n_343 & ~n_342) | (n_341 & n_342));
 assign n_182 = ((n_180 & ~n_179) | (n_178 & n_179));
 assign n_350 = ((n_348 & ~n_347) | (n_346 & n_347));
 assign n_177 = ((n_175 & ~n_174) | (n_173 & n_174));
 assign n_354 = ((n_353 & ~n_352) | (n_351 & n_352));
 assign n_172 = ((n_170 & ~n_467) | (n_168 & n_467));
 assign n_358 = ((n_357 & ~n_356) | (n_355 & n_356));
 assign n_167 = ((n_165 & ~n_164) | (n_163 & n_164));
 assign n_362 = ((n_361 & ~n_360) | (n_359 & n_360));
 assign n_162 = ((n_160 & ~n_159) | (n_158 & n_159));
 assign n_366 = ((n_365 & ~n_364) | (n_363 & n_364));
 assign n_157 = ((n_155 & ~n_154) | (n_153 & n_154));
 assign n_370 = ((n_369 & ~n_368) | (n_367 & n_368));
 assign n_152 = ((n_150 & ~n_149) | (n_148 & n_149));
 assign n_374 = ((n_373 & ~n_372) | (n_371 & n_372));
 assign n_147 = ((n_145 & ~n_144) | (n_143 & n_144));
 assign n_378 = ((n_377 & ~n_376) | (n_375 & n_376));
 assign n_142 = ((n_140 & ~n_466) | (n_138 & n_466));
 assign n_382 = ((n_381 & ~n_380) | (n_379 & n_380));
 assign n_137 = ((n_135 & ~n_134) | (n_133 & n_134));
 assign n_386 = ((n_385 & ~n_384) | (n_383 & n_384));
 assign n_132 = ((n_130 & ~n_129) | (n_128 & n_129));
 assign n_133 = ((n_131 & ~n_129) | ({in2[58]} & n_129));
 assign n_391 = ((n_389 & ~n_388) | (n_387 & n_388));
 assign n_127 = ((n_125 & ~n_465) | (n_123 & n_465));
 assign n_128 = ((n_126 & ~n_465) | ({in2[59]} & n_465));
 assign n_396 = ((n_394 & ~n_393) | (n_392 & n_393));
 assign n_122 = ((n_120 & ~n_464) | (n_450 & n_464));
 assign n_401 = ((n_399 & ~n_398) | (n_397 & n_398));
 assign {out1[14]} = ~n_342;
 assign {out1[1]} = ~n_398;
 assign {out1[2]} = ~n_393;
 assign {out1[3]} = ~n_388;
 assign {out1[4]} = ~n_384;
 assign {out1[5]} = ~n_380;
 assign {out1[6]} = ~n_376;
 assign {out1[7]} = ~n_372;
 assign {out1[8]} = ~n_368;
 assign {out1[9]} = ~n_364;
 assign {out1[10]} = ~n_360;
 assign {out1[11]} = ~n_356;
 assign {out1[12]} = ~n_352;
 assign {out1[13]} = ~n_347;
 assign {out1[30]} = ~n_268;
 assign {out1[16]} = ~n_334;
 assign {out1[17]} = ~n_330;
 assign {out1[18]} = ~n_326;
 assign {out1[19]} = ~n_322;
 assign n_117 = ((n_115 & ~n_463) | (n_451 & n_463));
 assign n_112 = ((n_110 & ~n_109) | (n_108 & n_109));
 assign sub_939_2_n_3 = (n_349 & n_452);
 assign sub_939_2_n_4 = ~(n_452 | n_349);
 assign sub_1546_2_n_4 = (n_35 | (n_402 & n_38));
 assign n_271 = ((n_269 & ~n_268) | (n_30 & n_268));
 assign sub_960_2_n_3 = (n_459 & n_344);
 assign sub_981_2_n_4 = ~(n_457 | n_46);
 assign n_47 = ((n_67 & ~stall) | (n_4 & stall));
 assign sub_1107_2_n_3 = (n_461 & n_40);
 assign sub_981_2_n_3 = (n_457 & n_46);
 assign sub_1107_2_n_4 = ~(n_461 | n_40);
 assign sub_1086_2_n_3 = (n_458 & n_41);
 assign sub_1086_2_n_4 = ~(n_458 | n_41);
 assign sub_1065_2_n_3 = (n_460 & n_42);
 assign sub_1065_2_n_4 = ~(n_460 | n_42);
 assign sub_1044_2_n_3 = (n_462 & n_43);
 assign sub_1023_2_n_3 = (n_455 & n_44);
 assign sub_1044_2_n_4 = ~(n_462 | n_43);
 assign sub_1023_2_n_4 = ~(n_455 | n_44);
 assign sub_1002_2_n_3 = (n_456 & n_45);
 assign sub_1002_2_n_4 = ~(n_456 | n_45);
 assign n_359 = ~(n_403 & (n_356 | sub_1317_2_n_2));
 assign n_333 = ~(n_404 & (n_330 | sub_1191_2_n_2));
 assign n_392 = ~(n_61 & (n_388 | sub_1485_2_n_2));
 assign n_341 = ~(n_405 & (n_338 | sub_1233_2_n_2));
 assign n_329 = ~(n_60 & (n_326 | sub_1170_2_n_2));
 assign n_367 = ~(n_62 & (n_364 | sub_1359_2_n_2));
 assign n_321 = ~(n_58 & (n_483 | sub_1128_2_n_2));
 assign n_387 = ~(n_395 & (n_384 | sub_1464_2_n_2));
 assign n_363 = ~(n_50 & (n_360 | sub_1338_2_n_2));
 assign sub_960_2_n_4 = ~(n_459 | n_344);
 assign n_325 = ~(n_390 & (n_322 | sub_1149_2_n_2));
 assign n_397 = ~(n_52 & (n_393 | sub_1506_2_n_2));
 assign n_337 = ~(n_53 & (n_334 | sub_1212_2_n_2));
 assign n_346 = ~(n_54 & (n_342 | sub_1254_2_n_2));
 assign n_375 = ~(n_55 & (n_372 | sub_1401_2_n_2));
 assign n_371 = ~(n_49 & (n_368 | sub_1380_2_n_2));
 assign n_351 = ~(n_56 & (n_347 | sub_1275_2_n_2));
 assign n_355 = ~(n_57 & (n_352 | sub_1296_2_n_2));
 assign n_383 = ~(n_59 & (n_380 | sub_1443_2_n_2));
 assign n_379 = ~(n_400 & (n_376 | sub_1422_2_n_2));
 assign n_402 = ~(n_63 & (n_398 | sub_1527_2_n_2));
 assign n_60 = ~(n_10 & (n_326 | n_51));
 assign n_63 = ~(n_2 & (n_398 | n_51));
 assign n_403 = ~(n_3 & (n_356 | n_51));
 assign n_404 = ~(n_5 & (n_330 | n_51));
 assign n_61 = ~(n_6 & (n_388 | n_51));
 assign n_405 = ~(n_8 & (n_338 | n_51));
 assign n_35 = (n_36 & n_4);
 assign n_62 = ~(n_11 & (n_364 | n_51));
 assign n_58 = ~(n_12 & (n_483 | n_51));
 assign n_395 = ~(n_13 & (n_384 | n_51));
 assign n_50 = ~(n_14 & (n_360 | n_51));
 assign n_390 = ~(n_20 & (n_322 | n_51));
 assign n_52 = ~(n_21 & (n_393 | n_51));
 assign n_53 = ~(n_22 & (n_334 | n_51));
 assign n_54 = ~(n_23 & (n_342 | n_51));
 assign n_55 = ~(n_24 & (n_372 | n_51));
 assign n_49 = ~(n_25 & (n_368 | n_51));
 assign n_56 = ~(n_26 & (n_347 | n_51));
 assign n_57 = ~(n_27 & (n_352 | n_51));
 assign n_59 = ~(n_28 & (n_380 | n_51));
 assign n_400 = ~(n_32 & (n_376 | n_51));
 assign n_34 = ~((n_68 & {in1[1]}) | (n_37 & stall));
 assign n_65 = ((n_265 & ~n_479) | (n_439 & n_479));
 assign n_268 = (n_267 ^ sub_918_2_n_9);
 assign sub_918_2_n_3 = ~(n_48 | ~n_30);
 assign sub_981_2_n_1 = ~(n_29 & n_51);
 assign sub_981_2_n_2 = ~(n_29 | n_51);
 assign sub_1107_2_n_1 = ~(n_51 & n_15);
 assign sub_1086_2_n_1 = ~(n_51 & n_17);
 assign sub_1065_2_n_2 = ~(n_51 | n_7);
 assign sub_939_2_n_2 = ~(n_9 | n_51);
 assign n_67 = ~({in1[0]} & ~{in2[0]});
 assign sub_960_2_n_2 = ~(n_31 | n_51);
 assign sub_1023_2_n_1 = ~(n_16 & n_51);
 assign sub_1086_2_n_2 = ~(n_51 | n_17);
 assign sub_1275_2_n_2 = (n_51 | n_26);
 assign sub_1128_2_n_2 = (n_51 | n_12);
 assign sub_1506_2_n_2 = (n_51 | n_21);
 assign sub_1254_2_n_2 = (n_51 | n_23);
 assign sub_1149_2_n_2 = (n_51 | n_20);
 assign sub_1233_2_n_2 = (n_51 | n_8);
 assign sub_1338_2_n_2 = (n_51 | n_14);
 assign sub_1401_2_n_2 = (n_51 | n_24);
 assign sub_1485_2_n_2 = (n_51 | n_6);
 assign sub_1212_2_n_2 = (n_51 | n_22);
 assign sub_1380_2_n_2 = (n_51 | n_25);
 assign sub_918_2_n_4 = ~(n_64 | n_30);
 assign sub_1002_2_n_2 = ~(n_18 | n_51);
 assign sub_1065_2_n_1 = ~(n_7 & n_51);
 assign sub_1044_2_n_1 = ~(n_19 & n_51);
 assign sub_1002_2_n_1 = ~(n_18 & n_51);
 assign sub_1044_2_n_2 = ~(n_19 | n_51);
 assign sub_918_2_n_2 = ~(n_51 | n_33);
 assign sub_939_2_n_1 = ~(n_9 & n_51);
 assign sub_1023_2_n_2 = ~(n_16 | n_51);
 assign sub_1107_2_n_2 = ~(n_51 | n_15);
 assign sub_918_2_n_1 = ~(n_51 & n_33);
 assign n_36 = ~(sub_1546_2_n_1 & n_39);
 assign sub_960_2_n_1 = ~(n_31 & n_51);
 assign sub_1443_2_n_2 = (n_51 | n_28);
 assign sub_1170_2_n_2 = (n_51 | n_10);
 assign sub_1422_2_n_2 = (n_51 | n_32);
 assign sub_1527_2_n_2 = (n_51 | n_2);
 assign sub_1317_2_n_2 = (n_51 | n_3);
 assign sub_1464_2_n_2 = (n_51 | n_13);
 assign sub_1359_2_n_2 = (n_51 | n_11);
 assign sub_1296_2_n_2 = (n_51 | n_27);
 assign sub_1191_2_n_2 = (n_51 | n_5);
 assign {out1[31]} = ~n_0;
 assign n_37 = ~n_38;
 assign n_38 = ~n_39;
 assign n_39 = ~sub_1527_2_n_1;
 assign sub_1527_2_n_1 = sub_1506_2_n_1;
 assign sub_1506_2_n_1 = sub_1485_2_n_1;
 assign sub_1485_2_n_1 = sub_1464_2_n_1;
 assign sub_1464_2_n_1 = sub_1443_2_n_1;
 assign sub_1443_2_n_1 = sub_1422_2_n_1;
 assign sub_1422_2_n_1 = sub_1401_2_n_1;
 assign sub_1401_2_n_1 = sub_1380_2_n_1;
 assign sub_1380_2_n_1 = sub_1359_2_n_1;
 assign sub_1359_2_n_1 = n_40;
 assign n_40 = sub_1338_2_n_1;
 assign sub_1338_2_n_1 = n_41;
 assign n_41 = n_42;
 assign n_42 = sub_1317_2_n_1;
 assign sub_1317_2_n_1 = n_43;
 assign n_43 = n_44;
 assign n_44 = sub_1296_2_n_1;
 assign sub_1296_2_n_1 = n_45;
 assign n_45 = n_46;
 assign n_46 = sub_1275_2_n_1;
 assign sub_1275_2_n_1 = n_344;
 assign n_344 = n_349;
 assign n_349 = sub_1254_2_n_1;
 assign sub_1254_2_n_1 = ~n_48;
 assign n_48 = ~n_64;
 assign n_64 = sub_1233_2_n_1;
 assign sub_1233_2_n_1 = sub_1212_2_n_1;
 assign sub_1212_2_n_1 = sub_1149_2_n_1;
 assign n_51 = ~n_1;
 assign n_68 = ~stall;
 assign n_106 = ~(sub_289_2_n_2 & ~{in1[1]});
 assign n_107 = ~((sub_289_2_n_1 & ~{in1[0]}) | ({in2[63]} & {in1[0]}));
 assign sub_289_2_n_2 = ~(sub_289_2_n_1 & {in1[0]});
 assign sub_289_2_n_1 = ~{in2[63]};
 assign n_109 = ~(sub_308_2_n_6 | sub_308_2_n_4);
 assign n_110 = ~(n_108 ^ ({in1[1]} ^ sub_308_2_n_3));
 assign sub_308_2_n_6 = ~(sub_308_2_n_2 | ~sub_308_2_n_3);
 assign n_111 = ~(sub_308_2_n_3 & ~(sub_308_2_n_0 & {in2[62]}));
 assign sub_308_2_n_4 = (sub_308_2_n_1 & n_108);
 assign sub_308_2_n_3 = ~({in1[0]} & ~{in2[62]});
 assign sub_308_2_n_2 = ~(n_108 | sub_308_2_n_1);
 assign sub_308_2_n_1 = ~{in1[1]};
 assign sub_308_2_n_0 = ~{in1[0]};
 assign sub_327_2_n_9 = ~(sub_327_2_n_4 | ~(sub_327_2_n_3 | sub_327_2_n_5));
 assign n_115 = ~(sub_327_2_n_7 ^ sub_327_2_n_3);
 assign sub_327_2_n_7 = ~(sub_327_2_n_4 | sub_327_2_n_5);
 assign n_116 = ~(sub_327_2_n_2 & ~sub_327_2_n_3);
 assign sub_327_2_n_5 = ~(n_451 | sub_327_2_n_1);
 assign sub_327_2_n_4 = (sub_327_2_n_1 & n_451);
 assign sub_327_2_n_3 = ~({in2[61]} | ~{in1[0]});
 assign sub_327_2_n_2 = ~({in2[61]} & ~{in1[0]});
 assign sub_327_2_n_1 = ~{in1[1]};
 assign sub_346_2_n_9 = ~(sub_346_2_n_7 | sub_346_2_n_3);
 assign n_120 = ~(sub_346_2_n_6 ^ sub_346_2_n_2);
 assign sub_346_2_n_7 = ~(sub_346_2_n_2 | sub_346_2_n_4);
 assign sub_346_2_n_6 = ~(sub_346_2_n_3 | sub_346_2_n_4);
 assign n_121 = ~(sub_346_2_n_1 & ~sub_346_2_n_2);
 assign sub_346_2_n_4 = ~(n_450 | ~{in1[1]});
 assign sub_346_2_n_3 = ~({in1[1]} | ~n_450);
 assign sub_346_2_n_2 = ~({in2[60]} | ~{in1[0]});
 assign sub_346_2_n_1 = ~({in2[60]} & ~{in1[0]});
 assign sub_365_2_n_5 = ((sub_365_2_n_3 & n_123) | ((n_123 & sub_365_2_n_2) | (sub_365_2_n_2 & sub_365_2_n_3)));
 assign n_125 = (n_123 ^ (sub_365_2_n_2 ^ sub_365_2_n_3));
 assign n_126 = ~(sub_365_2_n_3 & ~(sub_365_2_n_0 & {in2[59]}));
 assign sub_365_2_n_3 = ~({in1[0]} & ~{in2[59]});
 assign sub_365_2_n_2 = ~{in1[1]};
 assign sub_365_2_n_0 = ~{in1[0]};
 assign n_129 = ~(sub_384_2_n_4 ^ n_127);
 assign sub_384_2_n_4 = ((sub_384_2_n_2 & n_128) | ((n_128 & sub_384_2_n_1) | (sub_384_2_n_1 & sub_384_2_n_2)));
 assign n_130 = (n_128 ^ (sub_384_2_n_1 ^ sub_384_2_n_2));
 assign n_131 = ~(sub_384_2_n_2 & ~(sub_384_2_n_0 & {in2[58]}));
 assign sub_384_2_n_2 = ~({in1[0]} & ~{in2[58]});
 assign sub_384_2_n_1 = ~{in1[1]};
 assign sub_384_2_n_0 = ~{in1[0]};
 assign n_134 = ~(sub_403_2_n_4 ^ n_132);
 assign sub_403_2_n_4 = ((sub_403_2_n_2 & n_133) | ((n_133 & sub_403_2_n_1) | (sub_403_2_n_1 & sub_403_2_n_2)));
 assign n_135 = (n_133 ^ (sub_403_2_n_1 ^ sub_403_2_n_2));
 assign n_136 = ~(sub_403_2_n_2 & ~(sub_403_2_n_0 & {in2[57]}));
 assign sub_403_2_n_2 = ~({in1[0]} & ~{in2[57]});
 assign sub_403_2_n_1 = ~{in1[1]};
 assign sub_403_2_n_0 = ~{in1[0]};
 assign sub_422_2_n_5 = ((sub_422_2_n_3 & n_138) | ((n_138 & sub_422_2_n_2) | (sub_422_2_n_2 & sub_422_2_n_3)));
 assign n_140 = (n_138 ^ (sub_422_2_n_2 ^ sub_422_2_n_3));
 assign n_141 = ~(sub_422_2_n_3 & ~(sub_422_2_n_0 & {in2[56]}));
 assign sub_422_2_n_3 = ~({in1[0]} & ~{in2[56]});
 assign sub_422_2_n_2 = ~{in1[1]};
 assign sub_422_2_n_0 = ~{in1[0]};
 assign n_144 = ~(sub_441_2_n_4 ^ n_142);
 assign sub_441_2_n_4 = ((sub_441_2_n_2 & n_143) | ((n_143 & sub_441_2_n_1) | (sub_441_2_n_1 & sub_441_2_n_2)));
 assign n_145 = (n_143 ^ (sub_441_2_n_1 ^ sub_441_2_n_2));
 assign n_146 = ~(sub_441_2_n_2 & ~(sub_441_2_n_0 & {in2[55]}));
 assign sub_441_2_n_2 = ~({in1[0]} & ~{in2[55]});
 assign sub_441_2_n_1 = ~{in1[1]};
 assign sub_441_2_n_0 = ~{in1[0]};
 assign n_149 = ~(sub_460_2_n_4 ^ n_147);
 assign sub_460_2_n_4 = ((sub_460_2_n_2 & n_148) | ((n_148 & sub_460_2_n_1) | (sub_460_2_n_1 & sub_460_2_n_2)));
 assign n_150 = (n_148 ^ (sub_460_2_n_1 ^ sub_460_2_n_2));
 assign n_151 = ~(sub_460_2_n_2 & ~(sub_460_2_n_0 & {in2[54]}));
 assign sub_460_2_n_2 = ~({in1[0]} & ~{in2[54]});
 assign sub_460_2_n_1 = ~{in1[1]};
 assign sub_460_2_n_0 = ~{in1[0]};
 assign n_154 = ~(sub_479_2_n_6 & (sub_479_2_n_5 | n_152));
 assign sub_479_2_n_6 = ~(sub_479_2_n_5 & n_152);
 assign sub_479_2_n_5 = ((sub_479_2_n_2 & n_153) | ((n_153 & sub_479_2_n_1) | (sub_479_2_n_1 & sub_479_2_n_2)));
 assign n_155 = (n_153 ^ (sub_479_2_n_1 ^ sub_479_2_n_2));
 assign n_156 = ~(sub_479_2_n_2 & ~(sub_479_2_n_0 & {in2[53]}));
 assign sub_479_2_n_2 = ~({in1[0]} & ~{in2[53]});
 assign sub_479_2_n_1 = ~{in1[1]};
 assign sub_479_2_n_0 = ~{in1[0]};
 assign n_159 = ~(sub_498_2_n_4 ^ n_157);
 assign sub_498_2_n_4 = ((sub_498_2_n_2 & n_158) | ((n_158 & sub_498_2_n_1) | (sub_498_2_n_1 & sub_498_2_n_2)));
 assign n_160 = (n_158 ^ (sub_498_2_n_1 ^ sub_498_2_n_2));
 assign n_161 = ~(sub_498_2_n_2 & ~(sub_498_2_n_0 & {in2[52]}));
 assign sub_498_2_n_2 = ~({in1[0]} & ~{in2[52]});
 assign sub_498_2_n_1 = ~{in1[1]};
 assign sub_498_2_n_0 = ~{in1[0]};
 assign n_164 = ~(sub_517_2_n_4 ^ n_162);
 assign sub_517_2_n_4 = ((sub_517_2_n_2 & n_163) | ((n_163 & sub_517_2_n_1) | (sub_517_2_n_1 & sub_517_2_n_2)));
 assign n_165 = (n_163 ^ (sub_517_2_n_1 ^ sub_517_2_n_2));
 assign n_166 = ~(sub_517_2_n_2 & ~(sub_517_2_n_0 & {in2[51]}));
 assign sub_517_2_n_2 = ~({in1[0]} & ~{in2[51]});
 assign sub_517_2_n_1 = ~{in1[1]};
 assign sub_517_2_n_0 = ~{in1[0]};
 assign sub_536_2_n_5 = ((sub_536_2_n_3 & n_168) | ((n_168 & sub_536_2_n_2) | (sub_536_2_n_2 & sub_536_2_n_3)));
 assign n_170 = (n_168 ^ (sub_536_2_n_2 ^ sub_536_2_n_3));
 assign n_171 = ~(sub_536_2_n_3 & ~(sub_536_2_n_0 & {in2[50]}));
 assign sub_536_2_n_3 = ~({in1[0]} & ~{in2[50]});
 assign sub_536_2_n_2 = ~{in1[1]};
 assign sub_536_2_n_0 = ~{in1[0]};
 assign n_174 = ~(sub_555_2_n_4 ^ n_172);
 assign sub_555_2_n_4 = ((sub_555_2_n_2 & n_173) | ((n_173 & sub_555_2_n_1) | (sub_555_2_n_1 & sub_555_2_n_2)));
 assign n_175 = (n_173 ^ (sub_555_2_n_1 ^ sub_555_2_n_2));
 assign n_176 = ~(sub_555_2_n_2 & ~(sub_555_2_n_0 & {in2[49]}));
 assign sub_555_2_n_2 = ~({in1[0]} & ~{in2[49]});
 assign sub_555_2_n_1 = ~{in1[1]};
 assign sub_555_2_n_0 = ~{in1[0]};
 assign n_179 = ~(sub_574_2_n_4 ^ n_177);
 assign sub_574_2_n_4 = ((sub_574_2_n_2 & n_178) | ((n_178 & sub_574_2_n_1) | (sub_574_2_n_1 & sub_574_2_n_2)));
 assign n_180 = (n_178 ^ (sub_574_2_n_1 ^ sub_574_2_n_2));
 assign n_181 = ~(sub_574_2_n_2 & ~(sub_574_2_n_0 & {in2[48]}));
 assign sub_574_2_n_2 = ~({in1[0]} & ~{in2[48]});
 assign sub_574_2_n_1 = ~{in1[1]};
 assign sub_574_2_n_0 = ~{in1[0]};
 assign sub_593_2_n_5 = ((sub_593_2_n_3 & n_183) | ((n_183 & sub_593_2_n_2) | (sub_593_2_n_2 & sub_593_2_n_3)));
 assign n_185 = (n_183 ^ (sub_593_2_n_2 ^ sub_593_2_n_3));
 assign n_186 = ~(sub_593_2_n_3 & ~(sub_593_2_n_0 & {in2[47]}));
 assign sub_593_2_n_3 = ~({in1[0]} & ~{in2[47]});
 assign sub_593_2_n_2 = ~{in1[1]};
 assign sub_593_2_n_0 = ~{in1[0]};
 assign n_189 = ~(sub_612_2_n_4 ^ n_187);
 assign sub_612_2_n_4 = ((sub_612_2_n_2 & n_188) | ((n_188 & sub_612_2_n_1) | (sub_612_2_n_1 & sub_612_2_n_2)));
 assign n_190 = (n_188 ^ (sub_612_2_n_1 ^ sub_612_2_n_2));
 assign n_191 = ~(sub_612_2_n_2 & ~(sub_612_2_n_0 & {in2[46]}));
 assign sub_612_2_n_2 = ~({in1[0]} & ~{in2[46]});
 assign sub_612_2_n_1 = ~{in1[1]};
 assign sub_612_2_n_0 = ~{in1[0]};
 assign sub_631_2_n_5 = ((sub_631_2_n_3 & n_193) | ((n_193 & sub_631_2_n_2) | (sub_631_2_n_2 & sub_631_2_n_3)));
 assign n_195 = (n_193 ^ (sub_631_2_n_2 ^ sub_631_2_n_3));
 assign n_196 = ~(sub_631_2_n_3 & ~(sub_631_2_n_0 & {in2[45]}));
 assign sub_631_2_n_3 = ~({in1[0]} & ~{in2[45]});
 assign sub_631_2_n_2 = ~{in1[1]};
 assign sub_631_2_n_0 = ~{in1[0]};
 assign n_199 = ~(sub_650_2_n_4 ^ n_197);
 assign sub_650_2_n_4 = ((sub_650_2_n_2 & n_198) | ((n_198 & sub_650_2_n_1) | (sub_650_2_n_1 & sub_650_2_n_2)));
 assign n_200 = (n_198 ^ (sub_650_2_n_1 ^ sub_650_2_n_2));
 assign n_201 = ~(sub_650_2_n_2 & ~(sub_650_2_n_0 & {in2[44]}));
 assign sub_650_2_n_2 = ~({in1[0]} & ~{in2[44]});
 assign sub_650_2_n_1 = ~{in1[1]};
 assign sub_650_2_n_0 = ~{in1[0]};
 assign sub_669_2_n_5 = ((sub_669_2_n_3 & n_438) | ((n_438 & sub_669_2_n_2) | (sub_669_2_n_2 & sub_669_2_n_3)));
 assign n_205 = (n_438 ^ (sub_669_2_n_2 ^ sub_669_2_n_3));
 assign n_206 = ~(sub_669_2_n_3 & ~(sub_669_2_n_0 & {in2[43]}));
 assign sub_669_2_n_3 = ~({in1[0]} & ~{in2[43]});
 assign sub_669_2_n_2 = ~{in1[1]};
 assign sub_669_2_n_0 = ~{in1[0]};
 assign n_209 = (sub_688_2_n_8 ^ n_207);
 assign sub_688_2_n_8 = ~(sub_688_2_n_6 | sub_688_2_n_2);
 assign n_210 = ~(sub_688_2_n_5 ^ sub_688_2_n_1);
 assign sub_688_2_n_6 = ~(sub_688_2_n_1 | sub_688_2_n_3);
 assign sub_688_2_n_5 = ~(sub_688_2_n_2 | sub_688_2_n_3);
 assign n_211 = ~(sub_688_2_n_0 & ~sub_688_2_n_1);
 assign sub_688_2_n_3 = ~(n_208 | ~{in1[1]});
 assign sub_688_2_n_2 = ~({in1[1]} | ~n_208);
 assign sub_688_2_n_1 = ~({in2[42]} | ~{in1[0]});
 assign sub_688_2_n_0 = ~({in2[42]} & ~{in1[0]});
 assign sub_707_2_n_5 = ((sub_707_2_n_3 & n_437) | ((n_437 & sub_707_2_n_2) | (sub_707_2_n_2 & sub_707_2_n_3)));
 assign n_215 = (n_437 ^ (sub_707_2_n_2 ^ sub_707_2_n_3));
 assign n_216 = ~(sub_707_2_n_3 & ~(sub_707_2_n_0 & {in2[41]}));
 assign sub_707_2_n_3 = ~({in1[0]} & ~{in2[41]});
 assign sub_707_2_n_2 = ~{in1[1]};
 assign sub_707_2_n_0 = ~{in1[0]};
 assign n_219 = (sub_726_2_n_8 ^ n_217);
 assign sub_726_2_n_8 = ~(sub_726_2_n_6 | sub_726_2_n_2);
 assign n_220 = ~(sub_726_2_n_5 ^ sub_726_2_n_1);
 assign sub_726_2_n_6 = ~(sub_726_2_n_1 | sub_726_2_n_3);
 assign sub_726_2_n_5 = ~(sub_726_2_n_2 | sub_726_2_n_3);
 assign n_221 = ~(sub_726_2_n_0 & ~sub_726_2_n_1);
 assign sub_726_2_n_3 = ~(n_218 | ~{in1[1]});
 assign sub_726_2_n_2 = ~({in1[1]} | ~n_218);
 assign sub_726_2_n_1 = ~({in2[40]} | ~{in1[0]});
 assign sub_726_2_n_0 = ~({in2[40]} & ~{in1[0]});
 assign sub_745_2_n_5 = ((sub_745_2_n_3 & n_449) | ((n_449 & sub_745_2_n_2) | (sub_745_2_n_2 & sub_745_2_n_3)));
 assign n_225 = (n_449 ^ (sub_745_2_n_2 ^ sub_745_2_n_3));
 assign n_226 = ~(sub_745_2_n_3 & ~(sub_745_2_n_0 & {in2[39]}));
 assign sub_745_2_n_3 = ~({in1[0]} & ~{in2[39]});
 assign sub_745_2_n_2 = ~{in1[1]};
 assign sub_745_2_n_0 = ~{in1[0]};
 assign n_229 = (sub_764_2_n_8 ^ n_227);
 assign sub_764_2_n_8 = ~(sub_764_2_n_6 | sub_764_2_n_2);
 assign n_230 = ~(sub_764_2_n_5 ^ sub_764_2_n_1);
 assign sub_764_2_n_6 = ~(sub_764_2_n_1 | sub_764_2_n_3);
 assign sub_764_2_n_5 = ~(sub_764_2_n_2 | sub_764_2_n_3);
 assign n_231 = ~(sub_764_2_n_0 & ~sub_764_2_n_1);
 assign sub_764_2_n_3 = ~(n_448 | ~{in1[1]});
 assign sub_764_2_n_2 = ~({in1[1]} | ~n_448);
 assign sub_764_2_n_1 = ~({in2[38]} | ~{in1[0]});
 assign sub_764_2_n_0 = ~({in2[38]} & ~{in1[0]});
 assign sub_783_2_n_5 = ((sub_783_2_n_3 & n_446) | ((n_446 & sub_783_2_n_2) | (sub_783_2_n_2 & sub_783_2_n_3)));
 assign n_235 = (n_446 ^ (sub_783_2_n_2 ^ sub_783_2_n_3));
 assign n_236 = ~(sub_783_2_n_3 & ~(sub_783_2_n_0 & {in2[37]}));
 assign sub_783_2_n_3 = ~({in1[0]} & ~{in2[37]});
 assign sub_783_2_n_2 = ~{in1[1]};
 assign sub_783_2_n_0 = ~{in1[0]};
 assign sub_802_2_n_9 = ~(sub_802_2_n_7 | sub_802_2_n_3);
 assign n_240 = ~(sub_802_2_n_6 ^ sub_802_2_n_2);
 assign sub_802_2_n_7 = ~(sub_802_2_n_2 | sub_802_2_n_4);
 assign sub_802_2_n_6 = ~(sub_802_2_n_3 | sub_802_2_n_4);
 assign n_241 = ~(sub_802_2_n_1 & ~sub_802_2_n_2);
 assign sub_802_2_n_4 = ~(n_444 | ~{in1[1]});
 assign sub_802_2_n_3 = ~({in1[1]} | ~n_444);
 assign sub_802_2_n_2 = ~({in2[36]} | ~{in1[0]});
 assign sub_802_2_n_1 = ~({in2[36]} & ~{in1[0]});
 assign sub_821_2_n_9 = ~(sub_821_2_n_7 | sub_821_2_n_3);
 assign n_245 = ~(sub_821_2_n_6 ^ sub_821_2_n_2);
 assign sub_821_2_n_7 = ~(sub_821_2_n_2 | sub_821_2_n_4);
 assign sub_821_2_n_6 = ~(sub_821_2_n_3 | sub_821_2_n_4);
 assign n_246 = ~(sub_821_2_n_1 & ~sub_821_2_n_2);
 assign sub_821_2_n_4 = ~(n_443 | ~{in1[1]});
 assign sub_821_2_n_3 = ~({in1[1]} | ~n_443);
 assign sub_821_2_n_2 = ~({in2[35]} | ~{in1[0]});
 assign sub_821_2_n_1 = ~({in2[35]} & ~{in1[0]});
 assign sub_840_2_n_9 = ~(sub_840_2_n_7 | sub_840_2_n_3);
 assign n_250 = ~(sub_840_2_n_6 ^ sub_840_2_n_2);
 assign sub_840_2_n_7 = ~(sub_840_2_n_2 | sub_840_2_n_4);
 assign sub_840_2_n_6 = ~(sub_840_2_n_3 | sub_840_2_n_4);
 assign n_251 = ~(sub_840_2_n_1 & ~sub_840_2_n_2);
 assign sub_840_2_n_4 = ~(n_442 | ~{in1[1]});
 assign sub_840_2_n_3 = ~({in1[1]} | ~n_442);
 assign sub_840_2_n_2 = ~({in2[34]} | ~{in1[0]});
 assign sub_840_2_n_1 = ~({in2[34]} & ~{in1[0]});
 assign sub_859_2_n_9 = ~(sub_859_2_n_7 | sub_859_2_n_3);
 assign n_255 = ~(sub_859_2_n_6 ^ sub_859_2_n_2);
 assign sub_859_2_n_7 = ~(sub_859_2_n_2 | sub_859_2_n_4);
 assign sub_859_2_n_6 = ~(sub_859_2_n_3 | sub_859_2_n_4);
 assign n_256 = ~(sub_859_2_n_1 & ~sub_859_2_n_2);
 assign sub_859_2_n_4 = ~(n_441 | ~{in1[1]});
 assign sub_859_2_n_3 = ~({in1[1]} | ~n_441);
 assign sub_859_2_n_2 = ~({in2[33]} | ~{in1[0]});
 assign sub_859_2_n_1 = ~({in2[33]} & ~{in1[0]});
 assign sub_878_2_n_9 = ~(sub_878_2_n_7 | sub_878_2_n_3);
 assign n_260 = ~(sub_878_2_n_6 ^ sub_878_2_n_2);
 assign sub_878_2_n_7 = ~(sub_878_2_n_2 | sub_878_2_n_4);
 assign sub_878_2_n_6 = ~(sub_878_2_n_3 | sub_878_2_n_4);
 assign n_261 = ~(sub_878_2_n_1 & ~sub_878_2_n_2);
 assign sub_878_2_n_4 = ~(n_440 | ~{in1[1]});
 assign sub_878_2_n_3 = ~({in1[1]} | ~n_440);
 assign sub_878_2_n_2 = ~({in2[32]} | ~{in1[0]});
 assign sub_878_2_n_1 = ~({in2[32]} & ~{in1[0]});
 assign sub_897_2_n_9 = ~(sub_897_2_n_7 | sub_897_2_n_3);
 assign n_265 = ~(sub_897_2_n_6 ^ sub_897_2_n_2);
 assign sub_897_2_n_7 = ~(sub_897_2_n_2 | sub_897_2_n_4);
 assign sub_897_2_n_6 = ~(sub_897_2_n_3 | sub_897_2_n_4);
 assign n_266 = ~(sub_897_2_n_1 & ~sub_897_2_n_2);
 assign sub_897_2_n_4 = ~(n_439 | ~{in1[1]});
 assign sub_897_2_n_3 = ~({in1[1]} | ~n_439);
 assign sub_897_2_n_2 = ~({in2[31]} | ~{in1[0]});
 assign sub_897_2_n_1 = ~({in2[31]} & ~{in1[0]});
 assign sub_918_2_n_9 = ~(sub_918_2_n_7 | sub_918_2_n_3);
 assign n_269 = ~(sub_918_2_n_6 ^ sub_918_2_n_2);
 assign sub_918_2_n_7 = ~(sub_918_2_n_2 | sub_918_2_n_4);
 assign sub_918_2_n_6 = ~(sub_918_2_n_3 | sub_918_2_n_4);
 assign n_270 = ~(sub_918_2_n_1 & ~sub_918_2_n_2);
 assign sub_939_2_n_9 = ~(sub_939_2_n_7 | sub_939_2_n_3);
 assign n_274 = ~(sub_939_2_n_6 ^ sub_939_2_n_2);
 assign sub_939_2_n_7 = ~(sub_939_2_n_2 | sub_939_2_n_4);
 assign sub_939_2_n_6 = ~(sub_939_2_n_3 | sub_939_2_n_4);
 assign n_275 = ~(sub_939_2_n_1 & ~sub_939_2_n_2);
 assign sub_960_2_n_9 = ~(sub_960_2_n_7 | sub_960_2_n_3);
 assign n_279 = ~(sub_960_2_n_6 ^ sub_960_2_n_2);
 assign sub_960_2_n_7 = ~(sub_960_2_n_2 | sub_960_2_n_4);
 assign sub_960_2_n_6 = ~(sub_960_2_n_3 | sub_960_2_n_4);
 assign n_280 = ~(sub_960_2_n_1 & ~sub_960_2_n_2);
 assign n_283 = (sub_981_2_n_9 ^ n_281);
 assign sub_981_2_n_9 = ~(sub_981_2_n_7 | sub_981_2_n_3);
 assign n_284 = ~(sub_981_2_n_6 ^ sub_981_2_n_2);
 assign sub_981_2_n_7 = ~(sub_981_2_n_2 | sub_981_2_n_4);
 assign sub_981_2_n_6 = ~(sub_981_2_n_3 | sub_981_2_n_4);
 assign n_285 = ~(sub_981_2_n_1 & ~sub_981_2_n_2);
 assign n_288 = (sub_1002_2_n_9 ^ n_286);
 assign sub_1002_2_n_9 = ~(sub_1002_2_n_7 | sub_1002_2_n_3);
 assign n_289 = ~(sub_1002_2_n_6 ^ sub_1002_2_n_2);
 assign sub_1002_2_n_7 = ~(sub_1002_2_n_2 | sub_1002_2_n_4);
 assign sub_1002_2_n_6 = ~(sub_1002_2_n_3 | sub_1002_2_n_4);
 assign n_290 = ~(sub_1002_2_n_1 & ~sub_1002_2_n_2);
 assign n_293 = (sub_1023_2_n_9 ^ n_291);
 assign sub_1023_2_n_9 = ~(sub_1023_2_n_7 | sub_1023_2_n_3);
 assign n_294 = ~(sub_1023_2_n_6 ^ sub_1023_2_n_2);
 assign sub_1023_2_n_7 = ~(sub_1023_2_n_2 | sub_1023_2_n_4);
 assign sub_1023_2_n_6 = ~(sub_1023_2_n_3 | sub_1023_2_n_4);
 assign n_295 = ~(sub_1023_2_n_1 & ~sub_1023_2_n_2);
 assign n_298 = (sub_1044_2_n_9 ^ n_296);
 assign sub_1044_2_n_9 = ~(sub_1044_2_n_7 | sub_1044_2_n_3);
 assign n_299 = ~(sub_1044_2_n_6 ^ sub_1044_2_n_2);
 assign sub_1044_2_n_7 = ~(sub_1044_2_n_2 | sub_1044_2_n_4);
 assign sub_1044_2_n_6 = ~(sub_1044_2_n_3 | sub_1044_2_n_4);
 assign n_300 = ~(sub_1044_2_n_1 & ~sub_1044_2_n_2);
 assign n_303 = (sub_1065_2_n_9 ^ n_445);
 assign sub_1065_2_n_9 = ~(sub_1065_2_n_7 | sub_1065_2_n_3);
 assign n_304 = ~(sub_1065_2_n_6 ^ sub_1065_2_n_2);
 assign sub_1065_2_n_7 = ~(sub_1065_2_n_2 | sub_1065_2_n_4);
 assign sub_1065_2_n_6 = ~(sub_1065_2_n_3 | sub_1065_2_n_4);
 assign n_305 = ~(sub_1065_2_n_1 & ~sub_1065_2_n_2);
 assign n_308 = (sub_1086_2_n_9 ^ n_447);
 assign sub_1086_2_n_9 = ~(sub_1086_2_n_7 | sub_1086_2_n_3);
 assign n_309 = ~(sub_1086_2_n_6 ^ sub_1086_2_n_2);
 assign sub_1086_2_n_7 = ~(sub_1086_2_n_2 | sub_1086_2_n_4);
 assign sub_1086_2_n_6 = ~(sub_1086_2_n_3 | sub_1086_2_n_4);
 assign n_310 = ~(sub_1086_2_n_1 & ~sub_1086_2_n_2);
 assign n_313 = (sub_1107_2_n_9 ^ n_311);
 assign sub_1107_2_n_9 = ~(sub_1107_2_n_7 | sub_1107_2_n_3);
 assign n_314 = ~(sub_1107_2_n_6 ^ sub_1107_2_n_2);
 assign sub_1107_2_n_7 = ~(sub_1107_2_n_2 | sub_1107_2_n_4);
 assign sub_1107_2_n_6 = ~(sub_1107_2_n_3 | sub_1107_2_n_4);
 assign n_315 = ~(sub_1107_2_n_1 & ~sub_1107_2_n_2);
 assign sub_1128_2_n_5 = ((sub_1128_2_n_2 & n_453) | ((n_453 & sub_1149_2_n_1) | (sub_1149_2_n_1 & sub_1128_2_n_2)));
 assign n_319 = (n_453 ^ (sub_1149_2_n_1 ^ sub_1128_2_n_2));
 assign n_322 = ~(sub_1149_2_n_4 ^ n_320);
 assign sub_1149_2_n_4 = ((sub_1149_2_n_2 & n_321) | ((n_321 & sub_1149_2_n_1) | (sub_1149_2_n_1 & sub_1149_2_n_2)));
 assign n_323 = (n_321 ^ (sub_1149_2_n_1 ^ sub_1149_2_n_2));
 assign n_326 = ~(sub_1170_2_n_4 ^ n_324);
 assign sub_1170_2_n_4 = ((sub_1170_2_n_2 & n_325) | ((n_325 & sub_1149_2_n_1) | (sub_1149_2_n_1 & sub_1170_2_n_2)));
 assign n_327 = (n_325 ^ (sub_1149_2_n_1 ^ sub_1170_2_n_2));
 assign n_330 = ~(sub_1191_2_n_4 ^ n_328);
 assign sub_1191_2_n_4 = ((sub_1191_2_n_2 & n_329) | ((n_329 & sub_1149_2_n_1) | (sub_1149_2_n_1 & sub_1191_2_n_2)));
 assign n_331 = (n_329 ^ (sub_1149_2_n_1 ^ sub_1191_2_n_2));
 assign n_334 = ~(sub_1212_2_n_4 ^ n_332);
 assign sub_1212_2_n_4 = ((sub_1212_2_n_2 & n_333) | ((n_333 & sub_1212_2_n_1) | (sub_1212_2_n_1 & sub_1212_2_n_2)));
 assign n_335 = (n_333 ^ (sub_1212_2_n_1 ^ sub_1212_2_n_2));
 assign n_338 = ~(sub_1233_2_n_4 ^ n_336);
 assign sub_1233_2_n_4 = ((sub_1233_2_n_2 & n_337) | ((n_337 & sub_1233_2_n_1) | (sub_1233_2_n_1 & sub_1233_2_n_2)));
 assign n_339 = (n_337 ^ (sub_1233_2_n_1 ^ sub_1233_2_n_2));
 assign n_342 = ~(sub_1254_2_n_4 ^ n_340);
 assign sub_1254_2_n_4 = ((sub_1254_2_n_2 & n_341) | ((n_341 & sub_1254_2_n_1) | (sub_1254_2_n_1 & sub_1254_2_n_2)));
 assign n_343 = (n_341 ^ (sub_1254_2_n_1 ^ sub_1254_2_n_2));
 assign n_347 = ~(sub_1275_2_n_4 ^ n_345);
 assign sub_1275_2_n_4 = ((sub_1275_2_n_2 & n_346) | ((n_346 & sub_1275_2_n_1) | (sub_1275_2_n_1 & sub_1275_2_n_2)));
 assign n_348 = (n_346 ^ (sub_1275_2_n_1 ^ sub_1275_2_n_2));
 assign n_352 = ~(sub_1296_2_n_4 ^ n_350);
 assign sub_1296_2_n_4 = ((sub_1296_2_n_2 & n_351) | ((n_351 & sub_1296_2_n_1) | (sub_1296_2_n_1 & sub_1296_2_n_2)));
 assign n_353 = (n_351 ^ (sub_1296_2_n_1 ^ sub_1296_2_n_2));
 assign n_356 = ~(sub_1317_2_n_4 ^ n_354);
 assign sub_1317_2_n_4 = ((sub_1317_2_n_2 & n_355) | ((n_355 & sub_1317_2_n_1) | (sub_1317_2_n_1 & sub_1317_2_n_2)));
 assign n_357 = (n_355 ^ (sub_1317_2_n_1 ^ sub_1317_2_n_2));
 assign n_360 = ~(sub_1338_2_n_4 ^ n_358);
 assign sub_1338_2_n_4 = ((sub_1338_2_n_2 & n_359) | ((n_359 & sub_1338_2_n_1) | (sub_1338_2_n_1 & sub_1338_2_n_2)));
 assign n_361 = (n_359 ^ (sub_1338_2_n_1 ^ sub_1338_2_n_2));
 assign n_364 = ~(sub_1359_2_n_4 ^ n_362);
 assign sub_1359_2_n_4 = ((sub_1359_2_n_2 & n_363) | ((n_363 & sub_1359_2_n_1) | (sub_1359_2_n_1 & sub_1359_2_n_2)));
 assign n_365 = (n_363 ^ (sub_1359_2_n_1 ^ sub_1359_2_n_2));
 assign n_368 = ~(sub_1380_2_n_4 ^ n_366);
 assign sub_1380_2_n_4 = ((sub_1380_2_n_2 & n_367) | ((n_367 & sub_1380_2_n_1) | (sub_1380_2_n_1 & sub_1380_2_n_2)));
 assign n_369 = (n_367 ^ (sub_1380_2_n_1 ^ sub_1380_2_n_2));
 assign n_372 = ~(sub_1401_2_n_4 ^ n_370);
 assign sub_1401_2_n_4 = ((sub_1401_2_n_2 & n_371) | ((n_371 & sub_1401_2_n_1) | (sub_1401_2_n_1 & sub_1401_2_n_2)));
 assign n_373 = (n_371 ^ (sub_1401_2_n_1 ^ sub_1401_2_n_2));
 assign n_376 = ~(sub_1422_2_n_4 ^ n_374);
 assign sub_1422_2_n_4 = ((sub_1422_2_n_2 & n_375) | ((n_375 & sub_1422_2_n_1) | (sub_1422_2_n_1 & sub_1422_2_n_2)));
 assign n_377 = (n_375 ^ (sub_1422_2_n_1 ^ sub_1422_2_n_2));
 assign n_380 = ~(sub_1443_2_n_4 ^ n_378);
 assign sub_1443_2_n_4 = ((sub_1443_2_n_2 & n_379) | ((n_379 & sub_1443_2_n_1) | (sub_1443_2_n_1 & sub_1443_2_n_2)));
 assign n_381 = (n_379 ^ (sub_1443_2_n_1 ^ sub_1443_2_n_2));
 assign n_384 = ~(sub_1464_2_n_4 ^ n_382);
 assign sub_1464_2_n_4 = ((sub_1464_2_n_2 & n_383) | ((n_383 & sub_1464_2_n_1) | (sub_1464_2_n_1 & sub_1464_2_n_2)));
 assign n_385 = (n_383 ^ (sub_1464_2_n_1 ^ sub_1464_2_n_2));
 assign n_388 = ~(sub_1485_2_n_4 ^ n_386);
 assign sub_1485_2_n_4 = ((sub_1485_2_n_2 & n_387) | ((n_387 & sub_1485_2_n_1) | (sub_1485_2_n_1 & sub_1485_2_n_2)));
 assign n_389 = (n_387 ^ (sub_1485_2_n_1 ^ sub_1485_2_n_2));
 assign n_393 = ~(sub_1506_2_n_4 ^ n_391);
 assign sub_1506_2_n_4 = ((sub_1506_2_n_2 & n_392) | ((n_392 & sub_1506_2_n_1) | (sub_1506_2_n_1 & sub_1506_2_n_2)));
 assign n_394 = (n_392 ^ (sub_1506_2_n_1 ^ sub_1506_2_n_2));
 assign n_398 = ~(sub_1527_2_n_4 ^ n_396);
 assign sub_1527_2_n_4 = ((sub_1527_2_n_2 & n_397) | ((n_397 & sub_1527_2_n_1) | (sub_1527_2_n_1 & sub_1527_2_n_2)));
 assign n_399 = (n_397 ^ (sub_1527_2_n_1 ^ sub_1527_2_n_2));
 assign in2_190_2_ = ~(sub_1546_2_n_4 ^ n_401);
 assign sub_1546_2_n_1 = ~n_402;
 assign n_437 = ((n_211 & ~n_209) | ({in2[42]} & n_209));
 assign n_438 = ((n_201 & ~n_199) | ({in2[44]} & n_199));
 assign n_439 = ((n_261 & ~n_478) | ({in2[32]} & n_478));
 assign n_440 = ((n_256 & ~n_477) | ({in2[33]} & n_477));
 assign n_441 = ((n_251 & ~n_476) | ({in2[34]} & n_476));
 assign n_442 = ((n_246 & ~n_475) | ({in2[35]} & n_475));
 assign n_443 = ((n_241 & ~n_474) | ({in2[36]} & n_474));
 assign n_444 = ((n_236 & ~n_473) | ({in2[37]} & n_473));
 assign n_445 = ((n_299 & ~n_298) | (n_462 & n_298));
 assign n_446 = ((n_231 & ~n_229) | ({in2[38]} & n_229));
 assign n_447 = ((n_304 & ~n_303) | (n_460 & n_303));
 assign n_448 = ((n_226 & ~n_472) | ({in2[39]} & n_472));
 assign n_449 = ((n_221 & ~n_219) | ({in2[40]} & n_219));
 assign n_450 = ((n_116 & ~n_463) | ({in2[61]} & n_463));
 assign n_451 = ((n_111 & ~n_109) | ({in2[62]} & n_109));
 assign n_452 = ((n_270 & ~n_268) | (n_33 & n_268));
 assign n_453 = ((n_315 & ~n_313) | (n_15 & n_313));
 assign n_454 = ((n_266 & ~n_479) | ({in2[31]} & n_479));
 assign n_455 = ((n_290 & ~n_288) | (n_18 & n_288));
 assign n_456 = ((n_285 & ~n_283) | (n_29 & n_283));
 assign n_457 = ((n_280 & ~n_481) | (n_31 & n_481));
 assign n_458 = ((n_305 & ~n_303) | (n_7 & n_303));
 assign n_459 = ((n_275 & ~n_480) | (n_9 & n_480));
 assign n_460 = ((n_300 & ~n_298) | (n_19 & n_298));
 assign n_461 = ((n_310 & ~n_308) | (n_17 & n_308));
 assign n_462 = ((n_295 & ~n_293) | (n_16 & n_293));
 assign n_463 = (sub_327_2_n_9 ^ n_112);
 assign n_464 = (sub_346_2_n_9 ^ n_117);
 assign n_465 = ~(sub_365_2_n_5 ^ n_122);
 assign n_466 = ~(sub_422_2_n_5 ^ n_137);
 assign n_467 = ~(sub_536_2_n_5 ^ n_167);
 assign n_468 = ~(sub_593_2_n_5 ^ n_182);
 assign n_469 = ~(sub_631_2_n_5 ^ n_192);
 assign n_470 = ~(sub_669_2_n_5 ^ n_202);
 assign n_471 = ~(sub_707_2_n_5 ^ n_212);
 assign n_472 = ~(sub_745_2_n_5 ^ n_222);
 assign n_473 = ~(sub_783_2_n_5 ^ n_232);
 assign n_474 = (sub_802_2_n_9 ^ n_237);
 assign n_475 = (sub_821_2_n_9 ^ n_242);
 assign n_476 = (sub_840_2_n_9 ^ n_247);
 assign n_477 = (sub_859_2_n_9 ^ n_252);
 assign n_478 = (sub_878_2_n_9 ^ n_257);
 assign n_479 = (sub_897_2_n_9 ^ n_262);
 assign n_480 = (sub_939_2_n_9 ^ n_271);
 assign n_481 = (sub_960_2_n_9 ^ n_276);
 assign n_483 = (sub_1128_2_n_5 ^ n_482);
 assign n_482 = ~((n_314 & ~n_313) | (n_461 & n_313));
endmodule
