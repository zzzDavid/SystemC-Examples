`timescale 1ps / 1ps
module dut_entirecomputation_4(
          in1,
          in2,
          in3,
          in4,
          in5,
          in6,
          in7,
          in8,
          out1,
          clk,
          stall
);
   input [7:0] in1;
   input [7:0] in2;
   input [7:0] in3;
   input [7:0] in4;
   input [7:0] in5;
   input [7:0] in6;
   input [7:0] in7;
   input [7:0] in8;
   output [31:0] out1;
   input clk;
   input stall;
wire add_57_2_n_0, add_57_2_n_1, add_57_2_n_2, add_57_2_n_3, add_57_2_n_4,
     add_57_2_n_5, add_57_2_n_6, add_57_2_n_7, add_57_2_n_8, add_57_2_n_9,
     add_57_2_n_10, add_57_2_n_11, add_57_2_n_12, add_57_2_n_13, add_57_2_n_14,
     add_57_2_n_15, add_57_2_n_16, add_57_2_n_17, add_57_2_n_18, add_57_2_n_19,
     add_57_2_n_21, add_57_2_n_22, add_57_2_n_23, add_57_2_n_24, add_57_2_n_25,
     add_57_2_n_26, add_57_2_n_27, add_57_2_n_28, add_57_2_n_30, add_57_2_n_31,
     add_57_2_n_32, add_57_2_n_34, add_57_2_n_35, add_57_2_n_36, add_57_2_n_38,
     add_57_2_n_39, add_57_2_n_40, add_57_2_n_42, add_57_2_n_43, add_57_2_n_44,
     add_57_2_n_48, add_100_2_n_0, add_100_2_n_1, add_100_2_n_2, add_100_2_n_3,
     add_100_2_n_4, add_100_2_n_5, add_100_2_n_6, add_100_2_n_7, add_100_2_n_8,
     add_100_2_n_9, add_100_2_n_10, add_100_2_n_11, add_100_2_n_12,
     add_100_2_n_13, add_100_2_n_14, add_100_2_n_15, add_100_2_n_16,
     add_100_2_n_17, add_100_2_n_18, add_100_2_n_19, add_100_2_n_20,
     add_100_2_n_21, add_100_2_n_22, add_100_2_n_24, add_100_2_n_26,
     add_100_2_n_28, add_100_2_n_29, add_100_2_n_31, add_100_2_n_32,
     add_100_2_n_34, add_100_2_n_35, add_100_2_n_36, add_100_2_n_40,
     csa_tree_add_64_2_groupi_n_2, csa_tree_add_64_2_groupi_n_3,
     csa_tree_add_64_2_groupi_n_4, csa_tree_add_64_2_groupi_n_5,
     csa_tree_add_64_2_groupi_n_6, csa_tree_add_64_2_groupi_n_7,
     csa_tree_add_64_2_groupi_n_8, csa_tree_add_64_2_groupi_n_10,
     csa_tree_add_64_2_groupi_n_11, csa_tree_add_64_2_groupi_n_12,
     csa_tree_add_64_2_groupi_n_13, csa_tree_add_64_2_groupi_n_14,
     csa_tree_add_64_2_groupi_n_15, csa_tree_add_64_2_groupi_n_16,
     csa_tree_add_64_2_groupi_n_17, csa_tree_add_64_2_groupi_n_18,
     csa_tree_add_64_2_groupi_n_19, csa_tree_add_64_2_groupi_n_20,
     csa_tree_add_64_2_groupi_n_21, csa_tree_add_64_2_groupi_n_23,
     csa_tree_add_64_2_groupi_n_24, csa_tree_add_64_2_groupi_n_25,
     csa_tree_add_64_2_groupi_n_26, csa_tree_add_64_2_groupi_n_27,
     csa_tree_add_64_2_groupi_n_28, csa_tree_add_64_2_groupi_n_29,
     csa_tree_add_64_2_groupi_n_30, csa_tree_add_64_2_groupi_n_31,
     csa_tree_add_64_2_groupi_n_32, csa_tree_add_64_2_groupi_n_33,
     csa_tree_add_64_2_groupi_n_34, csa_tree_add_64_2_groupi_n_36,
     csa_tree_add_64_2_groupi_n_37, csa_tree_add_64_2_groupi_n_38,
     csa_tree_add_64_2_groupi_n_39, csa_tree_add_64_2_groupi_n_40,
     csa_tree_add_64_2_groupi_n_41, csa_tree_add_64_2_groupi_n_42,
     csa_tree_add_64_2_groupi_n_43, csa_tree_add_64_2_groupi_n_44,
     csa_tree_add_64_2_groupi_n_45, csa_tree_add_64_2_groupi_n_46,
     csa_tree_add_64_2_groupi_n_47, csa_tree_add_64_2_groupi_n_48,
     csa_tree_add_64_2_groupi_n_49, csa_tree_add_64_2_groupi_n_50,
     csa_tree_add_64_2_groupi_n_51, csa_tree_add_64_2_groupi_n_52,
     csa_tree_add_64_2_groupi_n_53, csa_tree_add_64_2_groupi_n_54,
     csa_tree_add_64_2_groupi_n_55, csa_tree_add_64_2_groupi_n_56,
     csa_tree_add_64_2_groupi_n_57, csa_tree_add_64_2_groupi_n_58,
     csa_tree_add_64_2_groupi_n_59, csa_tree_add_64_2_groupi_n_60,
     csa_tree_add_64_2_groupi_n_61, csa_tree_add_64_2_groupi_n_62,
     csa_tree_add_64_2_groupi_n_64, csa_tree_add_64_2_groupi_n_67,
     csa_tree_add_64_2_groupi_n_69, csa_tree_add_64_2_groupi_n_71,
     csa_tree_add_64_2_groupi_n_72, csa_tree_add_64_2_groupi_n_73,
     csa_tree_add_64_2_groupi_n_74, csa_tree_add_64_2_groupi_n_75,
     csa_tree_add_64_2_groupi_n_76, csa_tree_add_64_2_groupi_n_77,
     csa_tree_add_64_2_groupi_n_78, csa_tree_add_64_2_groupi_n_81,
     csa_tree_add_64_2_groupi_n_82, csa_tree_add_64_2_groupi_n_83,
     csa_tree_add_71_2_groupi_n_1, csa_tree_add_71_2_groupi_n_2,
     csa_tree_add_71_2_groupi_n_3, csa_tree_add_71_2_groupi_n_4,
     csa_tree_add_71_2_groupi_n_5, csa_tree_add_71_2_groupi_n_6,
     csa_tree_add_71_2_groupi_n_7, csa_tree_add_71_2_groupi_n_8,
     csa_tree_add_71_2_groupi_n_9, csa_tree_add_71_2_groupi_n_10,
     csa_tree_add_71_2_groupi_n_11, csa_tree_add_71_2_groupi_n_12,
     csa_tree_add_71_2_groupi_n_13, csa_tree_add_71_2_groupi_n_14,
     csa_tree_add_71_2_groupi_n_49, csa_tree_add_71_2_groupi_n_52,
     csa_tree_add_71_2_groupi_n_53, csa_tree_add_71_2_groupi_n_54,
     csa_tree_add_71_2_groupi_n_56, csa_tree_add_71_2_groupi_n_57,
     csa_tree_add_71_2_groupi_n_58, csa_tree_add_71_2_groupi_n_59,
     csa_tree_add_71_2_groupi_n_60, csa_tree_add_71_2_groupi_n_61,
     csa_tree_add_71_2_groupi_n_62, csa_tree_add_71_2_groupi_n_63,
     csa_tree_add_71_2_groupi_n_64, csa_tree_add_71_2_groupi_n_65,
     csa_tree_add_71_2_groupi_n_66, csa_tree_add_71_2_groupi_n_67,
     csa_tree_add_71_2_groupi_n_68, csa_tree_add_71_2_groupi_n_69,
     csa_tree_add_71_2_groupi_n_70, csa_tree_add_71_2_groupi_n_71,
     csa_tree_add_71_2_groupi_n_72, csa_tree_add_71_2_groupi_n_73,
     csa_tree_add_71_2_groupi_n_74, csa_tree_add_71_2_groupi_n_75,
     csa_tree_add_71_2_groupi_n_76, csa_tree_add_71_2_groupi_n_77,
     csa_tree_add_71_2_groupi_n_78, csa_tree_add_71_2_groupi_n_79,
     csa_tree_add_71_2_groupi_n_80, csa_tree_add_71_2_groupi_n_81,
     csa_tree_add_71_2_groupi_n_82, csa_tree_add_71_2_groupi_n_83,
     csa_tree_add_71_2_groupi_n_87, csa_tree_add_71_2_groupi_n_88,
     csa_tree_add_71_2_groupi_n_89, csa_tree_add_71_2_groupi_n_90,
     csa_tree_add_71_2_groupi_n_91, csa_tree_add_71_2_groupi_n_92,
     csa_tree_add_71_2_groupi_n_93, csa_tree_add_71_2_groupi_n_94,
     csa_tree_add_71_2_groupi_n_95, csa_tree_add_71_2_groupi_n_96,
     csa_tree_add_71_2_groupi_n_97, csa_tree_add_71_2_groupi_n_98,
     csa_tree_add_71_2_groupi_n_99, csa_tree_add_71_2_groupi_n_100,
     csa_tree_add_71_2_groupi_n_101, csa_tree_add_71_2_groupi_n_102,
     csa_tree_add_71_2_groupi_n_103, csa_tree_add_71_2_groupi_n_105,
     csa_tree_add_71_2_groupi_n_108, csa_tree_add_71_2_groupi_n_109,
     csa_tree_add_71_2_groupi_n_110, csa_tree_add_71_2_groupi_n_111,
     csa_tree_add_71_2_groupi_n_116, csa_tree_add_71_2_groupi_n_117,
     csa_tree_add_71_2_groupi_n_118, csa_tree_add_71_2_groupi_n_119,
     csa_tree_add_71_2_groupi_n_120, csa_tree_add_71_2_groupi_n_121,
     csa_tree_add_71_2_groupi_n_122, csa_tree_add_71_2_groupi_n_125,
     csa_tree_add_71_2_groupi_n_126, csa_tree_add_71_2_groupi_n_127,
     csa_tree_add_86_2_n_3, csa_tree_add_86_2_n_4, csa_tree_add_86_2_n_5,
     csa_tree_add_86_2_n_6, csa_tree_add_86_2_n_7, csa_tree_add_86_2_n_8,
     csa_tree_add_86_2_n_9, csa_tree_add_86_2_n_10, csa_tree_add_86_2_n_11,
     csa_tree_add_86_2_n_12, csa_tree_add_86_2_n_14, csa_tree_add_86_2_n_15,
     csa_tree_add_86_2_n_16, csa_tree_add_86_2_n_17, csa_tree_add_86_2_n_18,
     csa_tree_add_86_2_n_19, csa_tree_add_86_2_n_20, csa_tree_add_86_2_n_21,
     csa_tree_add_86_2_n_23, csa_tree_add_86_2_n_25, csa_tree_add_86_2_n_26,
     csa_tree_add_86_2_n_27, csa_tree_add_86_2_n_28, csa_tree_add_86_2_n_29,
     csa_tree_add_86_2_n_30, csa_tree_add_86_2_n_31, csa_tree_add_86_2_n_33,
     csa_tree_add_86_2_n_34, csa_tree_add_86_2_n_35, csa_tree_add_86_2_n_37,
     csa_tree_add_86_2_n_38, csa_tree_add_86_2_n_39, csa_tree_add_86_2_n_41,
     csa_tree_add_86_2_n_42, csa_tree_add_86_2_n_44, csa_tree_add_86_2_n_45,
     csa_tree_add_86_2_n_46, csa_tree_add_86_2_n_47, csa_tree_add_86_2_n_48,
     csa_tree_add_86_2_n_49, csa_tree_add_86_2_n_50, csa_tree_add_86_2_n_51,
     csa_tree_add_86_2_n_52, csa_tree_add_86_2_n_53, csa_tree_add_86_2_n_54,
     csa_tree_add_86_2_n_55, csa_tree_add_86_2_n_57, csa_tree_add_86_2_n_58,
     csa_tree_add_86_2_n_59, csa_tree_add_86_2_n_61, csa_tree_add_86_2_n_62,
     csa_tree_add_86_2_n_63, csa_tree_add_86_2_n_65, csa_tree_add_86_2_n_66,
     csa_tree_add_86_2_n_67, csa_tree_add_86_2_n_68, csa_tree_add_86_2_n_69,
     csa_tree_add_86_2_n_71, csa_tree_add_86_2_n_72, csa_tree_add_86_2_n_74,
     csa_tree_add_86_2_n_75, csa_tree_add_86_2_n_76, csa_tree_add_86_2_n_78,
     csa_tree_add_86_2_n_79, csa_tree_add_86_2_n_80, csa_tree_add_86_2_n_81,
     csa_tree_add_86_2_n_82, csa_tree_add_86_2_n_83, csa_tree_add_86_2_n_84,
     csa_tree_add_86_2_n_86, csa_tree_add_86_2_n_87, csa_tree_add_86_2_n_89,
     csa_tree_add_86_2_n_90, csa_tree_add_86_2_n_91, csa_tree_add_86_2_n_92,
     csa_tree_add_86_2_n_93, csa_tree_add_86_2_n_94, csa_tree_add_86_2_n_95,
     csa_tree_add_86_2_n_96, csa_tree_add_86_2_n_97, csa_tree_add_86_2_n_98,
     csa_tree_add_86_2_n_99, csa_tree_add_86_2_n_100, csa_tree_add_86_2_n_101,
     csa_tree_add_86_2_n_102, csa_tree_add_86_2_n_103, csa_tree_add_86_2_n_104,
     csa_tree_add_86_2_n_105, csa_tree_add_86_2_n_106, csa_tree_add_86_2_n_108,
     csa_tree_add_86_2_n_109, csa_tree_add_86_2_n_111, csa_tree_add_86_2_n_112,
     csa_tree_add_86_2_n_113, csa_tree_add_86_2_n_114, csa_tree_add_86_2_n_115,
     csa_tree_add_86_2_n_116, csa_tree_add_86_2_n_117, csa_tree_add_86_2_n_118,
     csa_tree_add_86_2_n_119, csa_tree_add_86_2_n_120, csa_tree_add_86_2_n_121,
     csa_tree_add_86_2_n_122, csa_tree_add_86_2_n_123, csa_tree_add_86_2_n_125,
     csa_tree_add_86_2_n_126, csa_tree_add_86_2_n_127, csa_tree_add_86_2_n_128,
     csa_tree_add_86_2_n_129, csa_tree_add_86_2_n_130, csa_tree_add_86_2_n_131,
     csa_tree_add_86_2_n_132, csa_tree_add_86_2_n_133, csa_tree_add_86_2_n_136,
     csa_tree_add_86_2_n_137, csa_tree_add_86_2_n_138, csa_tree_add_86_2_n_139,
     csa_tree_add_86_2_n_140, csa_tree_add_86_2_n_141, csa_tree_add_86_2_n_142,
     csa_tree_add_86_2_n_143, csa_tree_add_86_2_n_144, csa_tree_add_86_2_n_145,
     csa_tree_add_86_2_n_146, csa_tree_add_86_2_n_147, csa_tree_add_86_2_n_148,
     csa_tree_add_86_2_n_149, csa_tree_add_86_2_n_151, csa_tree_add_86_2_n_152,
     csa_tree_add_86_2_n_153, csa_tree_add_86_2_n_154, csa_tree_add_86_2_n_155,
     csa_tree_add_86_2_n_156, csa_tree_add_86_2_n_157, csa_tree_add_86_2_n_158,
     csa_tree_add_86_2_n_159, csa_tree_add_86_2_n_160, csa_tree_add_86_2_n_161,
     csa_tree_add_86_2_n_162, csa_tree_add_86_2_n_163, csa_tree_add_86_2_n_164,
     csa_tree_add_86_2_n_165, csa_tree_add_86_2_n_166, csa_tree_add_86_2_n_167,
     csa_tree_add_86_2_n_168, csa_tree_add_86_2_n_169, csa_tree_add_86_2_n_170,
     csa_tree_add_86_2_n_171, csa_tree_add_86_2_n_172, csa_tree_add_86_2_n_173,
     csa_tree_add_86_2_n_174, csa_tree_add_86_2_n_175, csa_tree_add_86_2_n_176,
     csa_tree_add_86_2_n_177, csa_tree_add_86_2_n_178, csa_tree_add_86_2_n_179,
     csa_tree_add_86_2_n_180, csa_tree_add_86_2_n_181, csa_tree_add_86_2_n_182,
     csa_tree_add_86_2_n_183, csa_tree_add_86_2_n_184, csa_tree_add_86_2_n_185,
     csa_tree_add_86_2_n_186, csa_tree_add_86_2_n_187, csa_tree_add_86_2_n_188,
     csa_tree_add_86_2_n_189, csa_tree_add_86_2_n_190, csa_tree_add_86_2_n_192,
     csa_tree_add_86_2_n_193, csa_tree_add_86_2_n_194, csa_tree_add_86_2_n_195,
     csa_tree_add_86_2_n_196, csa_tree_add_86_2_n_197, csa_tree_add_86_2_n_198,
     csa_tree_add_86_2_n_199, csa_tree_add_86_2_n_200, csa_tree_add_86_2_n_201,
     csa_tree_add_86_2_n_202, csa_tree_add_86_2_n_203, csa_tree_add_86_2_n_204,
     csa_tree_add_86_2_n_205, csa_tree_add_86_2_n_206, csa_tree_add_86_2_n_207,
     csa_tree_add_86_2_n_208, csa_tree_add_86_2_n_209, csa_tree_add_86_2_n_210,
     csa_tree_add_86_2_n_211, csa_tree_add_86_2_n_212, csa_tree_add_86_2_n_213,
     csa_tree_add_86_2_n_217, csa_tree_add_86_2_n_218, csa_tree_add_86_2_n_219,
     csa_tree_add_86_2_n_220, csa_tree_add_86_2_n_221, csa_tree_add_86_2_n_222,
     csa_tree_add_86_2_n_223, csa_tree_add_86_2_n_224, csa_tree_add_86_2_n_225,
     csa_tree_add_86_2_n_226, csa_tree_add_86_2_n_227, csa_tree_add_86_2_n_228,
     csa_tree_add_86_2_n_229, csa_tree_add_86_2_n_230, csa_tree_add_86_2_n_231,
     csa_tree_add_86_2_n_232, csa_tree_add_86_2_n_233, csa_tree_add_86_2_n_234,
     csa_tree_add_86_2_n_235, csa_tree_add_86_2_n_236, csa_tree_add_86_2_n_237,
     csa_tree_add_86_2_n_238, csa_tree_add_86_2_n_239, csa_tree_add_86_2_n_240,
     csa_tree_add_86_2_n_241, csa_tree_add_86_2_n_242, csa_tree_add_86_2_n_243,
     csa_tree_add_86_2_n_244, csa_tree_add_86_2_n_245, csa_tree_add_86_2_n_246,
     csa_tree_add_86_2_n_247, csa_tree_add_86_2_n_248, csa_tree_add_86_2_n_249,
     csa_tree_add_86_2_n_250, csa_tree_add_86_2_n_251, csa_tree_add_86_2_n_252,
     csa_tree_add_86_2_n_253, csa_tree_add_86_2_n_254, csa_tree_add_86_2_n_255,
     csa_tree_add_86_2_n_256, csa_tree_add_86_2_n_257, csa_tree_add_86_2_n_258,
     csa_tree_add_86_2_n_259, csa_tree_add_86_2_n_260, csa_tree_add_86_2_n_261,
     csa_tree_add_86_2_n_262, csa_tree_add_86_2_n_263, csa_tree_add_86_2_n_264,
     csa_tree_add_86_2_n_265, csa_tree_add_86_2_n_266, csa_tree_add_86_2_n_267,
     csa_tree_add_86_2_n_268, csa_tree_add_86_2_n_269, csa_tree_add_86_2_n_270,
     csa_tree_add_86_2_n_271, csa_tree_add_86_2_n_272, csa_tree_add_86_2_n_273,
     csa_tree_add_86_2_n_274, csa_tree_add_86_2_n_275, csa_tree_add_86_2_n_276,
     csa_tree_add_86_2_n_277, csa_tree_add_86_2_n_278, csa_tree_add_86_2_n_279,
     csa_tree_add_86_2_n_280, csa_tree_add_86_2_n_281, csa_tree_add_86_2_n_282,
     csa_tree_add_86_2_n_283, csa_tree_add_86_2_n_284, csa_tree_add_86_2_n_285,
     csa_tree_add_86_2_n_286, csa_tree_add_86_2_n_287, csa_tree_add_86_2_n_288,
     csa_tree_add_86_2_n_289, csa_tree_add_86_2_n_290, csa_tree_add_86_2_n_291,
     csa_tree_add_86_2_n_292, csa_tree_add_86_2_n_293, csa_tree_add_86_2_n_294,
     csa_tree_add_86_2_n_295, csa_tree_add_86_2_n_296, csa_tree_add_86_2_n_297,
     csa_tree_add_86_2_n_298, csa_tree_add_86_2_n_299, csa_tree_add_86_2_n_300,
     csa_tree_add_86_2_n_301, csa_tree_add_86_2_n_302, csa_tree_add_86_2_n_303,
     csa_tree_add_86_2_n_304, csa_tree_add_86_2_n_305, csa_tree_add_86_2_n_306,
     csa_tree_add_86_2_n_307, csa_tree_add_86_2_n_308, csa_tree_add_86_2_n_309,
     csa_tree_add_86_2_n_310, csa_tree_add_86_2_n_311, csa_tree_add_86_2_n_312,
     csa_tree_add_86_2_n_313, csa_tree_add_86_2_n_314, csa_tree_add_86_2_n_315,
     csa_tree_add_86_2_n_316, csa_tree_add_86_2_n_317, csa_tree_add_86_2_n_318,
     csa_tree_add_86_2_n_319, csa_tree_add_86_2_n_320, csa_tree_add_86_2_n_321,
     csa_tree_add_86_2_n_322, csa_tree_add_86_2_n_323, csa_tree_add_86_2_n_324,
     csa_tree_add_86_2_n_325, csa_tree_add_86_2_n_326, csa_tree_add_86_2_n_327,
     csa_tree_add_86_2_n_328, csa_tree_add_86_2_n_329, csa_tree_add_86_2_n_330,
     csa_tree_add_86_2_n_331, csa_tree_add_86_2_n_332, csa_tree_add_86_2_n_333,
     csa_tree_add_86_2_n_334, csa_tree_add_86_2_n_335, csa_tree_add_86_2_n_336,
     csa_tree_add_86_2_n_337, csa_tree_add_86_2_n_338, csa_tree_add_86_2_n_339,
     csa_tree_add_86_2_n_340, csa_tree_add_86_2_n_341, csa_tree_add_86_2_n_342,
     csa_tree_add_86_2_n_343, csa_tree_add_86_2_n_344, csa_tree_add_86_2_n_345,
     csa_tree_add_86_2_n_346, csa_tree_add_86_2_n_347, csa_tree_add_86_2_n_348,
     csa_tree_add_86_2_n_349, csa_tree_add_86_2_n_350, csa_tree_add_86_2_n_351,
     csa_tree_add_86_2_n_352, csa_tree_add_86_2_n_353, csa_tree_add_86_2_n_354,
     csa_tree_add_86_2_n_355, csa_tree_add_86_2_n_356, csa_tree_add_86_2_n_357,
     csa_tree_add_86_2_n_358, csa_tree_add_86_2_n_359, csa_tree_add_86_2_n_360,
     csa_tree_add_86_2_n_361, csa_tree_add_86_2_n_362, csa_tree_add_86_2_n_363,
     csa_tree_add_86_2_n_364, csa_tree_add_86_2_n_365, csa_tree_add_86_2_n_366,
     csa_tree_add_86_2_n_367, csa_tree_add_86_2_n_368, csa_tree_add_86_2_n_369,
     csa_tree_add_86_2_n_370, csa_tree_add_86_2_n_371, csa_tree_add_86_2_n_372,
     csa_tree_add_86_2_n_373, csa_tree_add_86_2_n_374, csa_tree_add_86_2_n_375,
     csa_tree_add_86_2_n_376, csa_tree_add_86_2_n_377, csa_tree_add_86_2_n_378,
     csa_tree_add_86_2_n_379, csa_tree_add_86_2_n_380, csa_tree_add_86_2_n_381,
     csa_tree_add_86_2_n_382, csa_tree_add_86_2_n_383, csa_tree_add_86_2_n_384,
     csa_tree_add_86_2_n_385, csa_tree_add_86_2_n_386, csa_tree_add_86_2_n_387,
     csa_tree_add_86_2_n_388, csa_tree_add_86_2_n_389, csa_tree_add_86_2_n_390,
     csa_tree_add_86_2_n_391, csa_tree_add_86_2_n_392, csa_tree_add_86_2_n_393,
     csa_tree_add_86_2_n_394, csa_tree_add_86_2_n_395, csa_tree_add_86_2_n_396,
     csa_tree_add_86_2_n_397, csa_tree_add_86_2_n_398, csa_tree_add_86_2_n_399,
     csa_tree_add_86_2_n_400, csa_tree_add_86_2_n_402, csa_tree_add_86_2_n_403,
     csa_tree_add_86_2_n_404, csa_tree_add_86_2_n_405, csa_tree_add_86_2_n_406,
     csa_tree_add_86_2_n_407, csa_tree_add_86_2_n_408, csa_tree_add_86_2_n_409,
     csa_tree_add_86_2_n_410, csa_tree_add_86_2_n_411, csa_tree_add_86_2_n_412,
     csa_tree_add_86_2_n_413, csa_tree_add_86_2_n_414, csa_tree_add_86_2_n_415,
     csa_tree_add_86_2_n_416, csa_tree_add_86_2_n_417, csa_tree_add_86_2_n_418,
     csa_tree_add_86_2_n_419, csa_tree_add_86_2_n_420, csa_tree_add_86_2_n_421,
     csa_tree_add_86_2_n_422, csa_tree_add_86_2_n_423, csa_tree_add_86_2_n_424,
     csa_tree_add_86_2_n_425, csa_tree_add_86_2_n_426, csa_tree_add_86_2_n_427,
     csa_tree_add_86_2_n_428, csa_tree_add_86_2_n_429, csa_tree_add_86_2_n_430,
     csa_tree_add_86_2_n_431, csa_tree_add_86_2_n_434, csa_tree_add_86_2_n_435,
     csa_tree_add_86_2_n_436, csa_tree_add_86_2_n_437, csa_tree_add_86_2_n_438,
     csa_tree_add_86_2_n_439, csa_tree_add_86_2_n_440, csa_tree_add_86_2_n_441,
     csa_tree_add_86_2_n_442, csa_tree_add_86_2_n_443, csa_tree_add_86_2_n_444,
     csa_tree_add_86_2_n_445, csa_tree_add_86_2_n_446, csa_tree_add_86_2_n_447,
     csa_tree_add_86_2_n_448, csa_tree_add_86_2_n_449, csa_tree_add_86_2_n_450,
     csa_tree_add_86_2_n_451, csa_tree_add_86_2_n_452, csa_tree_add_86_2_n_453,
     csa_tree_add_86_2_n_454, csa_tree_add_86_2_n_455, csa_tree_add_86_2_n_456,
     csa_tree_add_86_2_n_457, csa_tree_add_86_2_n_458, csa_tree_add_86_2_n_459,
     csa_tree_add_86_2_n_460, csa_tree_add_86_2_n_461, csa_tree_add_86_2_n_462,
     csa_tree_add_86_2_n_463, csa_tree_add_86_2_n_466, csa_tree_add_86_2_n_467,
     csa_tree_add_86_2_n_468, csa_tree_add_86_2_n_469, csa_tree_add_86_2_n_470,
     csa_tree_add_86_2_n_471, csa_tree_add_86_2_n_472, csa_tree_add_86_2_n_473,
     csa_tree_add_86_2_n_474, csa_tree_add_86_2_n_475, csa_tree_add_86_2_n_476,
     csa_tree_add_86_2_n_477, csa_tree_add_86_2_n_478, csa_tree_add_86_2_n_479,
     csa_tree_add_86_2_n_480, csa_tree_add_86_2_n_481, csa_tree_add_86_2_n_482,
     csa_tree_add_86_2_n_483, csa_tree_add_86_2_n_484, csa_tree_add_86_2_n_485,
     csa_tree_add_86_2_n_486, csa_tree_add_86_2_n_487, csa_tree_add_86_2_n_488,
     csa_tree_add_86_2_n_489, csa_tree_add_86_2_n_490, csa_tree_add_86_2_n_491,
     csa_tree_add_86_2_n_492, csa_tree_add_86_2_n_493, csa_tree_add_86_2_n_494,
     csa_tree_add_86_2_n_495, csa_tree_add_86_2_n_496, csa_tree_add_86_2_n_497,
     csa_tree_add_86_2_n_498, csa_tree_add_86_2_n_499, csa_tree_add_86_2_n_500,
     csa_tree_add_86_2_n_501, csa_tree_add_86_2_n_502, csa_tree_add_86_2_n_503,
     csa_tree_add_86_2_n_504, csa_tree_add_86_2_n_505, csa_tree_add_86_2_n_506,
     csa_tree_add_86_2_n_507, csa_tree_add_86_2_n_508, csa_tree_add_86_2_n_509,
     csa_tree_add_86_2_n_510, csa_tree_add_86_2_n_511, csa_tree_add_86_2_n_512,
     csa_tree_add_86_2_n_513, csa_tree_add_86_2_n_514, csa_tree_add_86_2_n_515,
     csa_tree_add_86_2_n_516, csa_tree_add_86_2_n_517, csa_tree_add_86_2_n_518,
     csa_tree_add_86_2_n_519, csa_tree_add_86_2_n_520, csa_tree_add_86_2_n_521,
     csa_tree_add_86_2_n_522, csa_tree_add_86_2_n_523, csa_tree_add_86_2_n_524,
     csa_tree_add_86_2_n_525, csa_tree_add_86_2_n_526, csa_tree_add_86_2_n_527,
     csa_tree_add_86_2_n_528, csa_tree_add_86_2_n_529, csa_tree_add_86_2_n_530,
     csa_tree_add_86_2_n_531, csa_tree_add_86_2_n_532, csa_tree_add_86_2_n_533,
     csa_tree_add_86_2_n_534, csa_tree_add_86_2_n_535, csa_tree_add_86_2_n_536,
     csa_tree_add_86_2_n_537, csa_tree_add_86_2_n_538, csa_tree_add_86_2_n_539,
     csa_tree_add_86_2_n_540, csa_tree_add_86_2_n_541, csa_tree_add_86_2_n_542,
     csa_tree_add_86_2_n_543, csa_tree_add_86_2_n_544, csa_tree_add_86_2_n_545,
     csa_tree_add_86_2_n_546, csa_tree_add_86_2_n_547, csa_tree_add_86_2_n_548,
     csa_tree_add_86_2_n_549, csa_tree_add_86_2_n_550, csa_tree_add_86_2_n_551,
     csa_tree_add_86_2_n_552, csa_tree_add_86_2_n_553, csa_tree_add_86_2_n_554,
     csa_tree_add_86_2_n_555, csa_tree_add_86_2_n_556, csa_tree_add_86_2_n_557,
     csa_tree_add_86_2_n_558, csa_tree_add_86_2_n_559, csa_tree_add_86_2_n_560,
     csa_tree_add_86_2_n_561, csa_tree_add_86_2_n_562, csa_tree_add_86_2_n_563,
     csa_tree_add_86_2_n_564, csa_tree_add_86_2_n_565, csa_tree_add_86_2_n_566,
     csa_tree_add_86_2_n_567, csa_tree_add_86_2_n_570, csa_tree_add_86_2_n_571,
     csa_tree_add_86_2_n_572, csa_tree_add_86_2_n_573, csa_tree_add_86_2_n_574,
     csa_tree_add_86_2_n_575, csa_tree_add_86_2_n_576, csa_tree_add_86_2_n_577,
     csa_tree_add_86_2_n_578, csa_tree_add_86_2_n_579, csa_tree_add_86_2_n_580,
     csa_tree_add_86_2_n_581, csa_tree_add_86_2_n_582, csa_tree_add_86_2_n_583,
     csa_tree_add_86_2_n_584, csa_tree_add_86_2_n_585, csa_tree_add_86_2_n_586,
     csa_tree_add_86_2_n_587, csa_tree_add_86_2_n_588, csa_tree_add_86_2_n_589,
     csa_tree_add_86_2_n_590, csa_tree_add_86_2_n_591, csa_tree_add_86_2_n_592,
     csa_tree_add_86_2_n_593, csa_tree_add_86_2_n_594, csa_tree_add_86_2_n_595,
     csa_tree_add_86_2_n_596, csa_tree_add_86_2_n_597, csa_tree_add_86_2_n_598,
     csa_tree_add_86_2_n_599, csa_tree_add_86_2_n_600, csa_tree_add_86_2_n_602,
     csa_tree_add_86_2_n_603, csa_tree_add_86_2_n_604, csa_tree_add_86_2_n_605,
     csa_tree_add_86_2_n_606, csa_tree_add_86_2_n_607, csa_tree_add_86_2_n_608,
     csa_tree_add_86_2_n_609, csa_tree_add_86_2_n_610, csa_tree_add_86_2_n_611,
     csa_tree_add_86_2_n_612, csa_tree_add_86_2_n_613, csa_tree_add_86_2_n_614,
     csa_tree_add_86_2_n_615, csa_tree_add_86_2_n_616, csa_tree_add_86_2_n_617,
     csa_tree_add_86_2_n_618, csa_tree_add_86_2_n_619, csa_tree_add_86_2_n_620,
     csa_tree_add_86_2_n_621, csa_tree_add_86_2_n_622, csa_tree_add_86_2_n_623,
     csa_tree_add_86_2_n_624, csa_tree_add_86_2_n_625, csa_tree_add_86_2_n_626,
     csa_tree_add_86_2_n_627, csa_tree_add_86_2_n_628, csa_tree_add_86_2_n_629,
     csa_tree_add_86_2_n_630, csa_tree_add_86_2_n_631, csa_tree_add_86_2_n_632,
     csa_tree_add_86_2_n_633, csa_tree_add_86_2_n_634, csa_tree_add_86_2_n_635,
     csa_tree_add_86_2_n_636, csa_tree_add_86_2_n_637, csa_tree_add_86_2_n_638,
     csa_tree_add_86_2_n_639, csa_tree_add_86_2_n_640, csa_tree_add_86_2_n_641,
     csa_tree_add_86_2_n_642, csa_tree_add_86_2_n_643, csa_tree_add_86_2_n_644,
     csa_tree_add_86_2_n_645, csa_tree_add_86_2_n_646, csa_tree_add_86_2_n_647,
     csa_tree_add_86_2_n_648, csa_tree_add_86_2_n_649, csa_tree_add_86_2_n_650,
     csa_tree_add_86_2_n_651, csa_tree_add_86_2_n_652, csa_tree_add_86_2_n_653,
     csa_tree_add_86_2_n_654, csa_tree_add_86_2_n_655, csa_tree_add_86_2_n_656,
     csa_tree_add_86_2_n_657, csa_tree_add_86_2_n_658, csa_tree_add_86_2_n_659,
     csa_tree_add_86_2_n_660, csa_tree_add_86_2_n_661, csa_tree_add_86_2_n_662,
     csa_tree_add_86_2_n_663, csa_tree_add_86_2_n_664, csa_tree_add_86_2_n_665,
     csa_tree_add_86_2_n_666, csa_tree_add_86_2_n_667, csa_tree_add_86_2_n_668,
     csa_tree_add_86_2_n_670, csa_tree_add_86_2_n_671, csa_tree_add_86_2_n_672,
     csa_tree_add_86_2_n_673, csa_tree_add_86_2_n_674, csa_tree_add_86_2_n_675,
     csa_tree_add_86_2_n_676, csa_tree_add_86_2_n_677, csa_tree_add_86_2_n_678,
     csa_tree_add_86_2_n_679, csa_tree_add_86_2_n_680, csa_tree_add_86_2_n_681,
     csa_tree_add_86_2_n_682, csa_tree_add_86_2_n_683, csa_tree_add_86_2_n_684,
     csa_tree_add_86_2_n_685, csa_tree_add_86_2_n_686, csa_tree_add_86_2_n_687,
     csa_tree_add_86_2_n_688, csa_tree_add_86_2_n_689, csa_tree_add_86_2_n_690,
     csa_tree_add_86_2_n_691, csa_tree_add_86_2_n_692, csa_tree_add_86_2_n_693,
     csa_tree_add_86_2_n_694, csa_tree_add_86_2_n_695, csa_tree_add_86_2_n_696,
     csa_tree_add_86_2_n_697, csa_tree_add_86_2_n_698, csa_tree_add_86_2_n_699,
     csa_tree_add_86_2_n_700, csa_tree_add_86_2_n_701, csa_tree_add_86_2_n_702,
     csa_tree_add_86_2_n_703, csa_tree_add_86_2_n_704, csa_tree_add_86_2_n_705,
     csa_tree_add_86_2_n_706, csa_tree_add_86_2_n_708, csa_tree_add_86_2_n_709,
     csa_tree_add_86_2_n_710, csa_tree_add_86_2_n_711, csa_tree_add_86_2_n_712,
     csa_tree_add_86_2_n_713, csa_tree_add_86_2_n_714, csa_tree_add_86_2_n_715,
     csa_tree_add_86_2_n_716, csa_tree_add_86_2_n_717, csa_tree_add_86_2_n_718,
     csa_tree_add_86_2_n_719, csa_tree_add_86_2_n_720, csa_tree_add_86_2_n_721,
     csa_tree_add_86_2_n_722, csa_tree_add_86_2_n_723, csa_tree_add_86_2_n_724,
     csa_tree_add_86_2_n_725, csa_tree_add_86_2_n_726, csa_tree_add_86_2_n_727,
     csa_tree_add_86_2_n_728, csa_tree_add_86_2_n_729, csa_tree_add_86_2_n_730,
     csa_tree_add_86_2_n_731, csa_tree_add_86_2_n_732, csa_tree_add_86_2_n_733,
     csa_tree_add_86_2_n_734, csa_tree_add_86_2_n_735, csa_tree_add_86_2_n_736,
     csa_tree_add_86_2_n_737, csa_tree_add_86_2_n_738, csa_tree_add_86_2_n_739,
     csa_tree_add_86_2_n_740, csa_tree_add_86_2_n_741, csa_tree_add_86_2_n_742,
     csa_tree_add_86_2_n_744, csa_tree_add_86_2_n_745, csa_tree_add_86_2_n_746,
     csa_tree_add_86_2_n_747, csa_tree_add_86_2_n_748, csa_tree_add_86_2_n_749,
     csa_tree_add_86_2_n_750, csa_tree_add_86_2_n_751, csa_tree_add_86_2_n_752,
     csa_tree_add_86_2_n_753, csa_tree_add_86_2_n_754, csa_tree_add_86_2_n_755,
     csa_tree_add_86_2_n_756, csa_tree_add_86_2_n_757, csa_tree_add_86_2_n_758,
     csa_tree_add_86_2_n_759, csa_tree_add_86_2_n_760, csa_tree_add_86_2_n_761,
     csa_tree_add_86_2_n_762, csa_tree_add_86_2_n_764, csa_tree_add_86_2_n_768,
     csa_tree_add_86_2_n_769, csa_tree_add_86_2_n_772, csa_tree_add_86_2_n_773,
     csa_tree_add_86_2_n_774, csa_tree_add_86_2_n_775, csa_tree_add_86_2_n_776,
     csa_tree_add_86_2_n_778, csa_tree_add_86_2_n_779, csa_tree_add_86_2_n_780,
     csa_tree_add_86_2_n_781, csa_tree_add_86_2_n_782, csa_tree_add_86_2_n_783,
     csa_tree_add_86_2_n_784, csa_tree_add_86_2_n_785, csa_tree_add_86_2_n_788,
     csa_tree_add_86_2_n_789, csa_tree_add_86_2_n_790, csa_tree_add_86_2_n_791,
     csa_tree_add_86_2_n_798, csa_tree_add_86_2_n_799, csa_tree_add_86_2_n_802,
     csa_tree_add_86_2_n_803, csa_tree_add_86_2_n_804, csa_tree_add_86_2_n_805,
     csa_tree_add_86_2_n_806, csa_tree_add_86_2_n_807, csa_tree_add_86_2_n_814,
     csa_tree_add_86_2_n_815, csa_tree_add_86_2_n_816, csa_tree_add_86_2_n_817,
     csa_tree_add_86_2_n_818, csa_tree_add_86_2_n_819, csa_tree_add_86_2_n_820,
     csa_tree_add_86_2_n_821, csa_tree_add_86_2_n_824, csa_tree_add_86_2_n_825,
     csa_tree_add_86_2_n_826, csa_tree_add_86_2_n_827, csa_tree_add_86_2_n_830,
     csa_tree_add_86_2_n_831, csa_tree_add_86_2_n_832, csa_tree_add_86_2_n_833,
     csa_tree_add_86_2_n_834, csa_tree_add_86_2_n_835, csa_tree_add_86_2_n_836,
     csa_tree_add_86_2_n_837, csa_tree_add_86_2_n_838, csa_tree_add_86_2_n_839,
     csa_tree_add_86_2_n_840, csa_tree_add_86_2_n_841, csa_tree_add_86_2_n_842,
     csa_tree_add_86_2_n_843, csa_tree_add_86_2_n_844, csa_tree_add_86_2_n_845,
     csa_tree_add_86_2_n_848, csa_tree_add_86_2_n_849, csa_tree_add_86_2_n_850,
     csa_tree_add_86_2_n_851, csa_tree_add_86_2_n_852, csa_tree_add_86_2_n_853,
     csa_tree_add_86_2_n_854, csa_tree_add_86_2_n_855, csa_tree_add_86_2_n_858,
     csa_tree_add_86_2_n_859, csa_tree_add_86_2_n_860, csa_tree_add_86_2_n_861,
     csa_tree_add_86_2_n_862, csa_tree_add_86_2_n_863, csa_tree_add_86_2_n_868,
     csa_tree_add_86_2_n_869, csa_tree_add_86_2_n_870, csa_tree_add_86_2_n_871,
     csa_tree_add_86_2_n_872, csa_tree_add_86_2_n_873, csa_tree_add_86_2_n_874,
     csa_tree_add_86_2_n_875, csa_tree_add_86_2_n_876, csa_tree_add_86_2_n_877,
     csa_tree_add_86_2_n_882, csa_tree_add_86_2_n_883, csa_tree_add_86_2_n_884,
     csa_tree_add_86_2_n_885, csa_tree_add_86_2_n_886, csa_tree_add_86_2_n_887,
     csa_tree_add_86_2_n_888, csa_tree_add_86_2_n_889, csa_tree_add_86_2_n_890,
     csa_tree_add_86_2_n_891, csa_tree_add_86_2_n_892, csa_tree_add_86_2_n_893,
     csa_tree_add_86_2_n_894, csa_tree_add_86_2_n_895, csa_tree_add_86_2_n_896,
     csa_tree_add_86_2_n_897, csa_tree_add_86_2_n_898, csa_tree_add_86_2_n_899,
     csa_tree_add_86_2_n_902, csa_tree_add_86_2_n_903, csa_tree_add_86_2_n_906,
     csa_tree_add_86_2_n_907, csa_tree_add_86_2_n_912, csa_tree_add_86_2_n_914,
     csa_tree_add_86_2_n_915, csa_tree_add_86_2_n_918, csa_tree_add_86_2_n_919,
     csa_tree_add_86_2_n_920, csa_tree_add_86_2_n_921, csa_tree_add_86_2_n_932,
     csa_tree_add_86_2_n_933, csa_tree_add_86_2_n_938, csa_tree_add_86_2_n_939,
     csa_tree_add_86_2_n_940, csa_tree_add_86_2_n_941, csa_tree_add_86_2_n_944,
     csa_tree_add_86_2_n_945, csa_tree_add_86_2_n_946, csa_tree_add_86_2_n_947,
     csa_tree_add_86_2_n_952, csa_tree_add_86_2_n_953, csa_tree_add_86_2_n_954,
     csa_tree_add_86_2_n_955, csa_tree_add_86_2_n_956, csa_tree_add_86_2_n_957,
     csa_tree_add_86_2_n_960, csa_tree_add_86_2_n_961, csa_tree_add_86_2_n_964,
     csa_tree_add_86_2_n_968, csa_tree_add_86_2_n_969, csa_tree_add_86_2_n_970,
     csa_tree_add_86_2_n_971, csa_tree_add_86_2_n_972, csa_tree_add_86_2_n_973,
     csa_tree_add_86_2_n_974, csa_tree_add_86_2_n_975, csa_tree_add_86_2_n_982,
     csa_tree_add_86_2_n_983, csa_tree_add_92_2_groupi_n_0,
     csa_tree_add_92_2_groupi_n_1, csa_tree_add_92_2_groupi_n_2,
     csa_tree_add_92_2_groupi_n_3, csa_tree_add_92_2_groupi_n_4,
     csa_tree_add_92_2_groupi_n_5, csa_tree_add_92_2_groupi_n_6,
     csa_tree_add_92_2_groupi_n_7, csa_tree_add_92_2_groupi_n_8,
     csa_tree_add_92_2_groupi_n_9, csa_tree_add_92_2_groupi_n_10,
     csa_tree_add_92_2_groupi_n_11, csa_tree_add_92_2_groupi_n_12,
     csa_tree_add_92_2_groupi_n_13, csa_tree_add_92_2_groupi_n_14,
     csa_tree_add_92_2_groupi_n_15, csa_tree_add_92_2_groupi_n_16,
     csa_tree_add_92_2_groupi_n_17, csa_tree_add_92_2_groupi_n_18,
     csa_tree_add_92_2_groupi_n_19, csa_tree_add_92_2_groupi_n_20,
     csa_tree_add_92_2_groupi_n_21, csa_tree_add_92_2_groupi_n_22,
     csa_tree_add_92_2_groupi_n_23, csa_tree_add_92_2_groupi_n_24,
     csa_tree_add_92_2_groupi_n_25, csa_tree_add_92_2_groupi_n_26,
     csa_tree_add_92_2_groupi_n_27, csa_tree_add_92_2_groupi_n_28,
     csa_tree_add_92_2_groupi_n_29, csa_tree_add_92_2_groupi_n_30,
     csa_tree_add_92_2_groupi_n_31, csa_tree_add_92_2_groupi_n_32,
     csa_tree_add_92_2_groupi_n_33, csa_tree_add_92_2_groupi_n_34,
     csa_tree_add_92_2_groupi_n_35, csa_tree_add_92_2_groupi_n_36,
     csa_tree_add_92_2_groupi_n_37, csa_tree_add_92_2_groupi_n_38,
     csa_tree_add_92_2_groupi_n_39, csa_tree_add_92_2_groupi_n_40,
     csa_tree_add_92_2_groupi_n_41, csa_tree_add_92_2_groupi_n_42,
     csa_tree_add_92_2_groupi_n_43, csa_tree_add_92_2_groupi_n_45,
     csa_tree_add_92_2_groupi_n_46, csa_tree_add_92_2_groupi_n_47,
     csa_tree_add_92_2_groupi_n_48, csa_tree_add_92_2_groupi_n_49,
     csa_tree_add_92_2_groupi_n_50, csa_tree_add_92_2_groupi_n_51,
     csa_tree_add_92_2_groupi_n_52, csa_tree_add_92_2_groupi_n_53,
     csa_tree_add_92_2_groupi_n_54, csa_tree_add_92_2_groupi_n_55,
     csa_tree_add_92_2_groupi_n_56, csa_tree_add_92_2_groupi_n_57,
     csa_tree_add_92_2_groupi_n_58, csa_tree_add_92_2_groupi_n_59,
     csa_tree_add_92_2_groupi_n_60, csa_tree_add_92_2_groupi_n_61,
     csa_tree_add_92_2_groupi_n_62, csa_tree_add_92_2_groupi_n_63,
     csa_tree_add_92_2_groupi_n_64, csa_tree_add_92_2_groupi_n_65,
     csa_tree_add_92_2_groupi_n_66, csa_tree_add_92_2_groupi_n_67,
     csa_tree_add_92_2_groupi_n_68, csa_tree_add_92_2_groupi_n_69,
     csa_tree_add_92_2_groupi_n_70, csa_tree_add_92_2_groupi_n_71,
     csa_tree_add_92_2_groupi_n_72, csa_tree_add_92_2_groupi_n_73,
     csa_tree_add_92_2_groupi_n_74, csa_tree_add_92_2_groupi_n_77,
     csa_tree_add_92_2_groupi_n_78, csa_tree_add_92_2_groupi_n_79,
     csa_tree_add_92_2_groupi_n_80, csa_tree_add_92_2_groupi_n_81,
     csa_tree_add_92_2_groupi_n_82, csa_tree_add_92_2_groupi_n_83,
     csa_tree_add_92_2_groupi_n_84, csa_tree_add_92_2_groupi_n_85,
     csa_tree_add_92_2_groupi_n_86, csa_tree_add_92_2_groupi_n_87,
     csa_tree_add_92_2_groupi_n_88, csa_tree_add_92_2_groupi_n_89,
     csa_tree_add_92_2_groupi_n_90, csa_tree_add_92_2_groupi_n_91,
     csa_tree_add_92_2_groupi_n_93, csa_tree_add_92_2_groupi_n_94,
     csa_tree_add_92_2_groupi_n_95, csa_tree_add_92_2_groupi_n_96,
     csa_tree_add_92_2_groupi_n_98, csa_tree_add_92_2_groupi_n_99,
     csa_tree_add_92_2_groupi_n_102, csa_tree_add_92_2_groupi_n_103,
     csa_tree_add_92_2_groupi_n_104, csa_tree_add_92_2_groupi_n_105,
     csa_tree_add_92_2_groupi_n_106, csa_tree_add_92_2_groupi_n_107,
     csa_tree_add_92_2_groupi_n_108, csa_tree_add_92_2_groupi_n_109,
     csa_tree_add_92_2_groupi_n_110, csa_tree_add_92_2_groupi_n_111,
     csa_tree_add_92_2_groupi_n_112, csa_tree_add_92_2_groupi_n_113,
     csa_tree_add_92_2_groupi_n_114, csa_tree_add_92_2_groupi_n_115,
     csa_tree_add_92_2_groupi_n_116, csa_tree_add_92_2_groupi_n_117,
     csa_tree_add_92_2_groupi_n_118, csa_tree_add_92_2_groupi_n_119,
     csa_tree_add_92_2_groupi_n_120, csa_tree_add_92_2_groupi_n_121,
     csa_tree_add_92_2_groupi_n_122, csa_tree_add_92_2_groupi_n_123,
     csa_tree_add_92_2_groupi_n_124, csa_tree_add_92_2_groupi_n_125,
     csa_tree_add_92_2_groupi_n_126, csa_tree_add_92_2_groupi_n_127,
     csa_tree_add_92_2_groupi_n_128, csa_tree_add_92_2_groupi_n_129,
     csa_tree_add_92_2_groupi_n_130, csa_tree_add_92_2_groupi_n_131,
     csa_tree_add_92_2_groupi_n_132, csa_tree_add_92_2_groupi_n_133,
     csa_tree_add_92_2_groupi_n_136, csa_tree_add_92_2_groupi_n_137,
     csa_tree_add_92_2_groupi_n_138, csa_tree_add_92_2_groupi_n_139,
     csa_tree_add_92_2_groupi_n_140, csa_tree_add_92_2_groupi_n_141,
     csa_tree_add_92_2_groupi_n_144, csa_tree_add_92_2_groupi_n_145,
     csa_tree_add_92_2_groupi_n_146, csa_tree_add_92_2_groupi_n_147,
     csa_tree_add_92_2_groupi_n_148, csa_tree_add_92_2_groupi_n_149,
     csa_tree_add_92_2_groupi_n_150, csa_tree_add_92_2_groupi_n_151,
     csa_tree_add_92_2_groupi_n_152, csa_tree_add_92_2_groupi_n_153,
     csa_tree_add_92_2_groupi_n_154, csa_tree_add_92_2_groupi_n_155,
     csa_tree_add_92_2_groupi_n_156, csa_tree_add_92_2_groupi_n_157,
     csa_tree_add_92_2_groupi_n_158, csa_tree_add_92_2_groupi_n_159,
     csa_tree_add_92_2_groupi_n_160, csa_tree_add_92_2_groupi_n_161,
     csa_tree_add_92_2_groupi_n_164, csa_tree_add_92_2_groupi_n_165,
     csa_tree_add_92_2_groupi_n_166, csa_tree_add_92_2_groupi_n_167,
     csa_tree_add_92_2_groupi_n_168, csa_tree_add_92_2_groupi_n_169,
     csa_tree_add_92_2_groupi_n_170, csa_tree_add_92_2_groupi_n_171,
     csa_tree_add_92_2_groupi_n_174, csa_tree_add_92_2_groupi_n_175,
     csa_tree_add_92_2_groupi_n_176, csa_tree_add_92_2_groupi_n_177,
     csa_tree_add_92_2_groupi_n_182, csa_tree_add_92_2_groupi_n_183,
     csa_tree_add_92_2_groupi_n_184, csa_tree_add_92_2_groupi_n_185,
     csa_tree_add_92_2_groupi_n_186, csa_tree_add_92_2_groupi_n_187,
     csa_tree_add_92_2_groupi_n_188, csa_tree_add_92_2_groupi_n_189,
     csa_tree_add_92_2_groupi_n_192, csa_tree_add_92_2_groupi_n_193,
     csa_tree_add_92_2_groupi_n_194, csa_tree_add_92_2_groupi_n_195,
     csa_tree_add_92_2_groupi_n_196, csa_tree_add_92_2_groupi_n_197,
     csa_tree_add_92_2_groupi_n_198, csa_tree_add_92_2_groupi_n_199,
     csa_tree_add_92_2_groupi_n_202, csa_tree_add_92_2_groupi_n_203,
     csa_tree_add_92_2_groupi_n_204, csa_tree_add_92_2_groupi_n_205,
     csa_tree_add_92_2_groupi_n_206, csa_tree_add_92_2_groupi_n_207,
     csa_tree_add_92_2_groupi_n_208, csa_tree_add_92_2_groupi_n_210,
     csa_tree_add_92_2_groupi_n_211, csa_tree_add_92_2_groupi_n_220,
     csa_tree_add_92_2_groupi_n_221, csa_tree_add_92_2_groupi_n_226,
     csa_tree_add_92_2_groupi_n_227, csa_tree_add_92_2_groupi_n_276,
     csa_tree_add_92_2_groupi_n_278, csa_tree_add_92_2_groupi_n_280,
     csa_tree_add_92_2_groupi_n_282, csa_tree_add_106_2_groupi_n_0,
     csa_tree_add_106_2_groupi_n_1, csa_tree_add_106_2_groupi_n_2,
     csa_tree_add_106_2_groupi_n_3, csa_tree_add_106_2_groupi_n_4,
     csa_tree_add_106_2_groupi_n_5, csa_tree_add_106_2_groupi_n_7,
     csa_tree_add_106_2_groupi_n_8, csa_tree_add_106_2_groupi_n_9,
     csa_tree_add_106_2_groupi_n_11, csa_tree_add_106_2_groupi_n_12,
     csa_tree_add_106_2_groupi_n_13, csa_tree_add_106_2_groupi_n_14,
     csa_tree_add_106_2_groupi_n_15, csa_tree_add_106_2_groupi_n_16,
     csa_tree_add_106_2_groupi_n_17, csa_tree_add_106_2_groupi_n_19,
     csa_tree_add_106_2_groupi_n_20, csa_tree_add_106_2_groupi_n_21,
     csa_tree_add_106_2_groupi_n_22, csa_tree_add_106_2_groupi_n_23,
     csa_tree_add_106_2_groupi_n_24, csa_tree_add_106_2_groupi_n_31,
     csa_tree_add_106_2_groupi_n_32, csa_tree_add_106_2_groupi_n_34,
     csa_tree_add_106_2_groupi_n_35, csa_tree_add_106_2_groupi_n_36,
     csa_tree_add_106_2_groupi_n_37, csa_tree_add_106_2_groupi_n_38,
     csa_tree_add_106_2_groupi_n_39, csa_tree_add_106_2_groupi_n_40,
     csa_tree_add_106_2_groupi_n_41, csa_tree_add_106_2_groupi_n_42,
     csa_tree_add_106_2_groupi_n_43, csa_tree_add_106_2_groupi_n_44,
     csa_tree_add_106_2_groupi_n_45, csa_tree_add_106_2_groupi_n_46,
     csa_tree_add_106_2_groupi_n_47, csa_tree_add_106_2_groupi_n_48,
     csa_tree_add_106_2_groupi_n_49, csa_tree_add_106_2_groupi_n_51,
     csa_tree_add_106_2_groupi_n_52, csa_tree_add_106_2_groupi_n_53,
     csa_tree_add_106_2_groupi_n_58, csa_tree_add_106_2_groupi_n_61,
     csa_tree_add_106_2_groupi_n_62, csa_tree_add_106_2_groupi_n_64,
     csa_tree_add_106_2_groupi_n_65, csa_tree_add_106_2_groupi_n_68,
     csa_tree_add_106_2_groupi_n_69, csa_tree_add_106_2_groupi_n_70,
     csa_tree_add_106_2_groupi_n_71, csa_tree_add_106_2_groupi_n_72,
     csa_tree_add_106_2_groupi_n_73, csa_tree_add_106_2_groupi_n_74,
     csa_tree_add_106_2_groupi_n_76, csa_tree_add_106_2_groupi_n_77,
     csa_tree_add_106_2_groupi_n_78, csa_tree_add_106_2_groupi_n_79,
     csa_tree_add_106_2_groupi_n_80, csa_tree_add_106_2_groupi_n_81,
     csa_tree_add_106_2_groupi_n_82, csa_tree_add_106_2_groupi_n_83,
     csa_tree_add_106_2_groupi_n_86, csa_tree_add_106_2_groupi_n_87,
     csa_tree_add_106_2_groupi_n_88, csa_tree_add_106_2_groupi_n_89,
     csa_tree_add_106_2_groupi_n_90, csa_tree_add_106_2_groupi_n_91,
     csa_tree_add_106_2_groupi_n_92, csa_tree_add_106_2_groupi_n_93,
     csa_tree_add_106_2_groupi_n_94, csa_tree_add_106_2_groupi_n_113,
     csa_tree_add_106_2_groupi_n_119, csa_tree_add_106_2_groupi_n_126,
     csa_tree_add_106_2_groupi_n_131, csa_tree_add_106_2_groupi_n_153,
     csa_tree_add_106_2_groupi_n_161, csa_tree_add_106_2_groupi_n_170,
     csa_tree_add_106_2_groupi_n_177, csa_tree_add_106_2_groupi_n_187,
     csa_tree_add_106_2_groupi_n_195, csa_tree_add_106_2_groupi_n_203,
     csa_tree_add_106_2_groupi_n_207, csa_tree_add_106_2_groupi_n_208,
     csa_tree_add_106_2_groupi_n_211, csa_tree_add_106_2_groupi_n_212,
     csa_tree_add_106_2_groupi_n_215, csa_tree_add_106_2_groupi_n_217,
     csa_tree_add_106_2_groupi_n_218, csa_tree_add_106_2_groupi_n_220,
     csa_tree_add_106_2_groupi_n_221, csa_tree_add_106_2_groupi_n_222,
     csa_tree_add_106_2_groupi_n_223, csa_tree_add_106_2_groupi_n_224,
     csa_tree_add_106_2_groupi_n_225, csa_tree_add_106_2_groupi_n_226,
     csa_tree_add_106_2_groupi_n_227, csa_tree_add_106_2_groupi_n_228,
     csa_tree_add_106_2_groupi_n_229, csa_tree_add_106_2_groupi_n_230,
     csa_tree_add_106_2_groupi_n_233, csa_tree_add_106_2_groupi_n_240,
     csa_tree_add_106_2_groupi_n_245, csa_tree_add_106_2_groupi_n_248,
     csa_tree_add_106_2_groupi_n_262, csa_tree_add_106_2_groupi_n_268,
     csa_tree_add_106_2_groupi_n_311, csa_tree_add_106_2_groupi_n_312,
     csa_tree_add_106_2_groupi_n_332, csa_tree_add_106_2_groupi_n_333,
     csa_tree_add_106_2_groupi_n_335, csa_tree_add_106_2_groupi_n_336,
     csa_tree_add_106_2_groupi_n_337, csa_tree_add_106_2_groupi_n_338,
     csa_tree_add_106_2_groupi_n_343, csa_tree_add_106_2_groupi_n_344,
     csa_tree_add_106_2_groupi_n_345, csa_tree_add_106_2_groupi_n_346,
     csa_tree_add_106_2_groupi_n_347, csa_tree_add_106_2_groupi_n_348,
     csa_tree_add_106_2_groupi_n_349, csa_tree_add_106_2_groupi_n_350,
     csa_tree_add_106_2_groupi_n_353, csa_tree_add_106_2_groupi_n_362,
     csa_tree_add_106_2_groupi_n_364, csa_tree_add_106_2_groupi_n_365,
     csa_tree_add_106_2_groupi_n_366, csa_tree_add_106_2_groupi_n_367,
     csa_tree_add_106_2_groupi_n_368, csa_tree_add_106_2_groupi_n_369,
     csa_tree_add_106_2_groupi_n_370, csa_tree_add_106_2_groupi_n_371,
     csa_tree_add_106_2_groupi_n_372, csa_tree_add_106_2_groupi_n_373,
     csa_tree_add_106_2_groupi_n_374, csa_tree_add_106_2_groupi_n_375,
     csa_tree_add_106_2_groupi_n_376, csa_tree_add_106_2_groupi_n_377,
     csa_tree_add_106_2_groupi_n_378, csa_tree_add_106_2_groupi_n_380,
     csa_tree_add_106_2_groupi_n_381, csa_tree_add_106_2_groupi_n_382,
     csa_tree_add_106_2_groupi_n_383, csa_tree_add_106_2_groupi_n_384,
     csa_tree_add_106_2_groupi_n_385, csa_tree_add_106_2_groupi_n_386,
     csa_tree_add_106_2_groupi_n_387, csa_tree_add_106_2_groupi_n_389,
     csa_tree_add_106_2_groupi_n_390, csa_tree_add_106_2_groupi_n_391,
     csa_tree_add_106_2_groupi_n_392, csa_tree_add_106_2_groupi_n_393,
     csa_tree_add_106_2_groupi_n_394, csa_tree_add_106_2_groupi_n_395,
     csa_tree_add_106_2_groupi_n_397, csa_tree_add_106_2_groupi_n_398,
     csa_tree_add_106_2_groupi_n_399, csa_tree_add_106_2_groupi_n_401,
     csa_tree_add_106_2_groupi_n_402, csa_tree_add_106_2_groupi_n_403,
     csa_tree_add_106_2_groupi_n_404, csa_tree_add_106_2_groupi_n_405,
     csa_tree_add_106_2_groupi_n_408, csa_tree_add_106_2_groupi_n_409,
     csa_tree_add_106_2_groupi_n_411, csa_tree_add_106_2_groupi_n_412,
     csa_tree_add_106_2_groupi_n_413, csa_tree_add_106_2_groupi_n_414,
     csa_tree_add_106_2_groupi_n_415, csa_tree_add_106_2_groupi_n_416,
     csa_tree_add_106_2_groupi_n_417, csa_tree_add_106_2_groupi_n_418,
     csa_tree_add_106_2_groupi_n_420, csa_tree_add_106_2_groupi_n_421,
     csa_tree_add_106_2_groupi_n_422, csa_tree_add_106_2_groupi_n_423,
     csa_tree_add_106_2_groupi_n_424, csa_tree_add_106_2_groupi_n_425,
     csa_tree_add_106_2_groupi_n_426, csa_tree_add_106_2_groupi_n_427,
     csa_tree_add_106_2_groupi_n_428, csa_tree_add_106_2_groupi_n_429,
     csa_tree_add_106_2_groupi_n_430, csa_tree_add_106_2_groupi_n_431,
     csa_tree_add_106_2_groupi_n_432, csa_tree_add_106_2_groupi_n_433,
     csa_tree_add_106_2_groupi_n_434, csa_tree_add_106_2_groupi_n_435,
     csa_tree_add_106_2_groupi_n_436, csa_tree_add_106_2_groupi_n_437,
     csa_tree_add_106_2_groupi_n_440, csa_tree_add_106_2_groupi_n_441,
     csa_tree_add_106_2_groupi_n_442, csa_tree_add_106_2_groupi_n_443,
     csa_tree_add_106_2_groupi_n_446, csa_tree_add_106_2_groupi_n_447,
     csa_tree_add_106_2_groupi_n_448, csa_tree_add_106_2_groupi_n_449,
     csa_tree_add_106_2_groupi_n_450, csa_tree_add_106_2_groupi_n_451,
     csa_tree_add_106_2_groupi_n_452, csa_tree_add_106_2_groupi_n_453,
     csa_tree_add_106_2_groupi_n_454, csa_tree_add_106_2_groupi_n_455,
     csa_tree_add_106_2_groupi_n_457, csa_tree_add_106_2_groupi_n_458,
     csa_tree_add_106_2_groupi_n_460, csa_tree_add_106_2_groupi_n_461,
     csa_tree_add_106_2_groupi_n_462, csa_tree_add_106_2_groupi_n_463,
     csa_tree_add_106_2_groupi_n_464, csa_tree_add_106_2_groupi_n_465,
     csa_tree_add_106_2_groupi_n_467, csa_tree_add_106_2_groupi_n_468,
     csa_tree_add_106_2_groupi_n_470, csa_tree_add_106_2_groupi_n_471,
     csa_tree_add_106_2_groupi_n_472, csa_tree_add_106_2_groupi_n_475,
     csa_tree_add_106_2_groupi_n_476, csa_tree_add_106_2_groupi_n_477,
     csa_tree_add_106_2_groupi_n_478, csa_tree_add_106_2_groupi_n_479,
     csa_tree_add_106_2_groupi_n_480, csa_tree_add_106_2_groupi_n_481,
     csa_tree_add_106_2_groupi_n_482, csa_tree_add_106_2_groupi_n_483,
     csa_tree_add_106_2_groupi_n_484, csa_tree_add_106_2_groupi_n_485,
     csa_tree_add_106_2_groupi_n_486, csa_tree_add_106_2_groupi_n_488,
     csa_tree_add_106_2_groupi_n_489, csa_tree_add_106_2_groupi_n_490,
     csa_tree_add_106_2_groupi_n_491, csa_tree_add_106_2_groupi_n_492,
     csa_tree_add_106_2_groupi_n_494, csa_tree_add_106_2_groupi_n_495,
     csa_tree_add_106_2_groupi_n_496, csa_tree_add_106_2_groupi_n_497,
     csa_tree_add_106_2_groupi_n_499, csa_tree_add_106_2_groupi_n_500,
     csa_tree_add_106_2_groupi_n_501, csa_tree_add_106_2_groupi_n_502,
     csa_tree_add_106_2_groupi_n_503, csa_tree_add_106_2_groupi_n_504,
     csa_tree_add_106_2_groupi_n_506, csa_tree_add_106_2_groupi_n_507,
     csa_tree_add_106_2_groupi_n_508, csa_tree_add_106_2_groupi_n_510,
     csa_tree_add_106_2_groupi_n_511, csa_tree_add_106_2_groupi_n_512,
     csa_tree_add_106_2_groupi_n_513, csa_tree_add_106_2_groupi_n_514,
     csa_tree_add_106_2_groupi_n_515, csa_tree_add_106_2_groupi_n_516,
     csa_tree_add_106_2_groupi_n_517, csa_tree_add_106_2_groupi_n_520,
     csa_tree_add_106_2_groupi_n_521, csa_tree_add_106_2_groupi_n_523,
     csa_tree_add_106_2_groupi_n_524, csa_tree_add_106_2_groupi_n_526,
     csa_tree_add_106_2_groupi_n_527, csa_tree_add_106_2_groupi_n_528,
     csa_tree_add_106_2_groupi_n_529, csa_tree_add_106_2_groupi_n_530,
     csa_tree_add_106_2_groupi_n_531, csa_tree_add_106_2_groupi_n_532,
     csa_tree_add_106_2_groupi_n_533, csa_tree_add_106_2_groupi_n_534,
     csa_tree_add_106_2_groupi_n_535, csa_tree_add_106_2_groupi_n_536,
     csa_tree_add_106_2_groupi_n_538, csa_tree_add_106_2_groupi_n_539,
     csa_tree_add_106_2_groupi_n_540, csa_tree_add_106_2_groupi_n_542,
     csa_tree_add_106_2_groupi_n_543, csa_tree_add_106_2_groupi_n_544,
     csa_tree_add_106_2_groupi_n_546, csa_tree_add_106_2_groupi_n_547,
     csa_tree_add_106_2_groupi_n_549, csa_tree_add_106_2_groupi_n_550,
     csa_tree_add_106_2_groupi_n_551, csa_tree_add_106_2_groupi_n_553,
     csa_tree_add_106_2_groupi_n_554, csa_tree_add_106_2_groupi_n_555,
     csa_tree_add_106_2_groupi_n_556, csa_tree_add_106_2_groupi_n_558,
     csa_tree_add_106_2_groupi_n_559, csa_tree_add_106_2_groupi_n_562,
     csa_tree_add_106_2_groupi_n_563, csa_tree_add_106_2_groupi_n_564,
     csa_tree_add_106_2_groupi_n_565, csa_tree_add_106_2_groupi_n_566,
     csa_tree_add_106_2_groupi_n_567, csa_tree_add_106_2_groupi_n_568,
     csa_tree_add_106_2_groupi_n_569, csa_tree_add_106_2_groupi_n_570,
     csa_tree_add_106_2_groupi_n_571, csa_tree_add_106_2_groupi_n_572,
     csa_tree_add_106_2_groupi_n_573, csa_tree_add_106_2_groupi_n_574,
     csa_tree_add_106_2_groupi_n_575, csa_tree_add_106_2_groupi_n_577,
     csa_tree_add_106_2_groupi_n_578, csa_tree_add_106_2_groupi_n_579,
     csa_tree_add_106_2_groupi_n_581, csa_tree_add_106_2_groupi_n_582,
     csa_tree_add_106_2_groupi_n_583, csa_tree_add_106_2_groupi_n_584,
     csa_tree_add_106_2_groupi_n_585, csa_tree_add_106_2_groupi_n_586,
     csa_tree_add_106_2_groupi_n_587, csa_tree_add_106_2_groupi_n_588,
     csa_tree_add_106_2_groupi_n_589, csa_tree_add_106_2_groupi_n_590,
     csa_tree_add_106_2_groupi_n_592, csa_tree_add_106_2_groupi_n_596,
     csa_tree_add_106_2_groupi_n_598, csa_tree_add_106_2_groupi_n_599,
     csa_tree_add_106_2_groupi_n_600, csa_tree_add_106_2_groupi_n_601,
     csa_tree_add_106_2_groupi_n_602, csa_tree_add_106_2_groupi_n_603,
     csa_tree_add_106_2_groupi_n_604, csa_tree_add_106_2_groupi_n_605,
     csa_tree_add_106_2_groupi_n_606, csa_tree_add_106_2_groupi_n_607,
     csa_tree_add_106_2_groupi_n_608, csa_tree_add_106_2_groupi_n_609,
     csa_tree_add_106_2_groupi_n_610, csa_tree_add_106_2_groupi_n_612,
     csa_tree_add_106_2_groupi_n_613, csa_tree_add_106_2_groupi_n_614,
     csa_tree_add_106_2_groupi_n_615, csa_tree_add_106_2_groupi_n_616,
     csa_tree_add_106_2_groupi_n_617, csa_tree_add_106_2_groupi_n_618,
     csa_tree_add_106_2_groupi_n_619, csa_tree_add_106_2_groupi_n_620,
     csa_tree_add_106_2_groupi_n_621, csa_tree_add_106_2_groupi_n_622,
     csa_tree_add_106_2_groupi_n_623, csa_tree_add_106_2_groupi_n_624,
     csa_tree_add_106_2_groupi_n_625, csa_tree_add_106_2_groupi_n_626,
     csa_tree_add_106_2_groupi_n_628, csa_tree_add_106_2_groupi_n_630,
     csa_tree_add_106_2_groupi_n_631, csa_tree_add_106_2_groupi_n_632,
     csa_tree_add_106_2_groupi_n_633, csa_tree_add_106_2_groupi_n_634,
     csa_tree_add_106_2_groupi_n_635, csa_tree_add_106_2_groupi_n_636,
     csa_tree_add_106_2_groupi_n_637, csa_tree_add_106_2_groupi_n_638,
     csa_tree_add_106_2_groupi_n_639, csa_tree_add_106_2_groupi_n_640,
     csa_tree_add_106_2_groupi_n_641, csa_tree_add_106_2_groupi_n_642,
     csa_tree_add_106_2_groupi_n_643, csa_tree_add_106_2_groupi_n_644,
     csa_tree_add_106_2_groupi_n_645, csa_tree_add_106_2_groupi_n_646,
     csa_tree_add_106_2_groupi_n_647, csa_tree_add_106_2_groupi_n_648,
     csa_tree_add_106_2_groupi_n_649, csa_tree_add_106_2_groupi_n_650,
     csa_tree_add_106_2_groupi_n_651, csa_tree_add_106_2_groupi_n_652,
     csa_tree_add_106_2_groupi_n_653, csa_tree_add_106_2_groupi_n_654,
     csa_tree_add_106_2_groupi_n_655, csa_tree_add_106_2_groupi_n_656,
     csa_tree_add_106_2_groupi_n_657, csa_tree_add_106_2_groupi_n_658,
     csa_tree_add_106_2_groupi_n_659, csa_tree_add_106_2_groupi_n_660,
     csa_tree_add_106_2_groupi_n_661, csa_tree_add_106_2_groupi_n_662,
     csa_tree_add_106_2_groupi_n_663, csa_tree_add_106_2_groupi_n_664,
     csa_tree_add_106_2_groupi_n_665, csa_tree_add_106_2_groupi_n_666,
     csa_tree_add_106_2_groupi_n_667, csa_tree_add_106_2_groupi_n_668,
     csa_tree_add_106_2_groupi_n_669, csa_tree_add_106_2_groupi_n_670,
     csa_tree_add_106_2_groupi_n_671, csa_tree_add_106_2_groupi_n_672,
     csa_tree_add_106_2_groupi_n_673, csa_tree_add_106_2_groupi_n_674,
     csa_tree_add_106_2_groupi_n_675, csa_tree_add_106_2_groupi_n_676,
     csa_tree_add_106_2_groupi_n_677, csa_tree_add_106_2_groupi_n_678,
     csa_tree_add_106_2_groupi_n_679, csa_tree_add_106_2_groupi_n_680,
     csa_tree_add_106_2_groupi_n_681, csa_tree_add_106_2_groupi_n_682,
     csa_tree_add_106_2_groupi_n_683, csa_tree_add_106_2_groupi_n_684,
     csa_tree_add_106_2_groupi_n_685, csa_tree_add_106_2_groupi_n_686,
     csa_tree_add_106_2_groupi_n_687, csa_tree_add_106_2_groupi_n_688,
     csa_tree_add_106_2_groupi_n_689, csa_tree_add_106_2_groupi_n_690,
     csa_tree_add_106_2_groupi_n_691, csa_tree_add_106_2_groupi_n_693,
     csa_tree_add_106_2_groupi_n_696, csa_tree_add_106_2_groupi_n_697,
     csa_tree_add_106_2_groupi_n_698, csa_tree_add_106_2_groupi_n_699,
     csa_tree_add_106_2_groupi_n_700, csa_tree_add_106_2_groupi_n_701,
     csa_tree_add_106_2_groupi_n_702, csa_tree_add_106_2_groupi_n_703,
     csa_tree_add_106_2_groupi_n_704, csa_tree_add_106_2_groupi_n_705,
     csa_tree_add_106_2_groupi_n_706, csa_tree_add_106_2_groupi_n_707,
     csa_tree_add_106_2_groupi_n_708, csa_tree_add_106_2_groupi_n_709,
     csa_tree_add_106_2_groupi_n_710, csa_tree_add_106_2_groupi_n_711,
     csa_tree_add_106_2_groupi_n_712, csa_tree_add_106_2_groupi_n_713,
     csa_tree_add_106_2_groupi_n_714, csa_tree_add_106_2_groupi_n_715,
     csa_tree_add_106_2_groupi_n_716, csa_tree_add_106_2_groupi_n_717,
     csa_tree_add_106_2_groupi_n_718, csa_tree_add_106_2_groupi_n_719,
     csa_tree_add_106_2_groupi_n_720, csa_tree_add_106_2_groupi_n_721,
     csa_tree_add_106_2_groupi_n_722, csa_tree_add_106_2_groupi_n_723,
     csa_tree_add_106_2_groupi_n_724, csa_tree_add_106_2_groupi_n_727,
     csa_tree_add_106_2_groupi_n_728, csa_tree_add_106_2_groupi_n_729,
     csa_tree_add_106_2_groupi_n_730, csa_tree_add_106_2_groupi_n_731,
     csa_tree_add_106_2_groupi_n_732, csa_tree_add_106_2_groupi_n_733,
     csa_tree_add_106_2_groupi_n_734, csa_tree_add_106_2_groupi_n_735,
     csa_tree_add_106_2_groupi_n_736, csa_tree_add_106_2_groupi_n_737,
     csa_tree_add_106_2_groupi_n_738, csa_tree_add_106_2_groupi_n_739,
     csa_tree_add_106_2_groupi_n_740, csa_tree_add_106_2_groupi_n_741,
     csa_tree_add_106_2_groupi_n_742, csa_tree_add_106_2_groupi_n_743,
     csa_tree_add_106_2_groupi_n_744, csa_tree_add_106_2_groupi_n_745,
     csa_tree_add_106_2_groupi_n_746, csa_tree_add_106_2_groupi_n_747,
     csa_tree_add_106_2_groupi_n_748, csa_tree_add_106_2_groupi_n_749,
     csa_tree_add_106_2_groupi_n_750, csa_tree_add_106_2_groupi_n_751,
     csa_tree_add_106_2_groupi_n_752, csa_tree_add_106_2_groupi_n_753,
     csa_tree_add_106_2_groupi_n_754, csa_tree_add_106_2_groupi_n_757,
     csa_tree_add_106_2_groupi_n_758, csa_tree_add_106_2_groupi_n_761,
     csa_tree_add_106_2_groupi_n_762, csa_tree_add_106_2_groupi_n_763,
     csa_tree_add_106_2_groupi_n_764, csa_tree_add_106_2_groupi_n_767,
     csa_tree_add_106_2_groupi_n_768, csa_tree_add_106_2_groupi_n_769,
     csa_tree_add_106_2_groupi_n_770, csa_tree_add_106_2_groupi_n_771,
     csa_tree_add_106_2_groupi_n_772, csa_tree_add_106_2_groupi_n_773,
     csa_tree_add_106_2_groupi_n_774, csa_tree_add_106_2_groupi_n_775,
     csa_tree_add_106_2_groupi_n_776, csa_tree_add_106_2_groupi_n_777,
     csa_tree_add_106_2_groupi_n_778, csa_tree_add_106_2_groupi_n_779,
     csa_tree_add_106_2_groupi_n_780, csa_tree_add_106_2_groupi_n_781,
     csa_tree_add_106_2_groupi_n_782, csa_tree_add_106_2_groupi_n_783,
     csa_tree_add_106_2_groupi_n_784, csa_tree_add_106_2_groupi_n_785,
     csa_tree_add_106_2_groupi_n_786, csa_tree_add_106_2_groupi_n_787,
     csa_tree_add_106_2_groupi_n_788, csa_tree_add_106_2_groupi_n_789,
     csa_tree_add_106_2_groupi_n_791, csa_tree_add_106_2_groupi_n_792,
     csa_tree_add_106_2_groupi_n_795, csa_tree_add_106_2_groupi_n_796,
     csa_tree_add_106_2_groupi_n_797, csa_tree_add_106_2_groupi_n_798,
     csa_tree_add_106_2_groupi_n_801, csa_tree_add_106_2_groupi_n_802,
     csa_tree_add_106_2_groupi_n_805, csa_tree_add_106_2_groupi_n_806,
     csa_tree_add_106_2_groupi_n_807, csa_tree_add_106_2_groupi_n_808,
     csa_tree_add_106_2_groupi_n_809, csa_tree_add_106_2_groupi_n_810,
     csa_tree_add_106_2_groupi_n_811, csa_tree_add_106_2_groupi_n_812,
     csa_tree_add_106_2_groupi_n_813, csa_tree_add_106_2_groupi_n_814,
     csa_tree_add_106_2_groupi_n_815, csa_tree_add_106_2_groupi_n_816,
     csa_tree_add_106_2_groupi_n_817, csa_tree_add_106_2_groupi_n_818,
     csa_tree_add_106_2_groupi_n_819, csa_tree_add_106_2_groupi_n_820,
     csa_tree_add_106_2_groupi_n_821, csa_tree_add_106_2_groupi_n_822,
     csa_tree_add_106_2_groupi_n_823, csa_tree_add_106_2_groupi_n_824,
     csa_tree_add_106_2_groupi_n_825, csa_tree_add_106_2_groupi_n_830,
     csa_tree_add_106_2_groupi_n_832, csa_tree_add_106_2_groupi_n_833,
     csa_tree_add_106_2_groupi_n_834, csa_tree_add_106_2_groupi_n_835,
     csa_tree_add_106_2_groupi_n_838, csa_tree_add_106_2_groupi_n_839,
     csa_tree_add_106_2_groupi_n_840, csa_tree_add_106_2_groupi_n_841,
     csa_tree_add_106_2_groupi_n_842, csa_tree_add_106_2_groupi_n_843,
     csa_tree_add_106_2_groupi_n_844, csa_tree_add_106_2_groupi_n_845,
     csa_tree_add_106_2_groupi_n_850, csa_tree_add_106_2_groupi_n_851,
     csa_tree_add_106_2_groupi_n_852, csa_tree_add_106_2_groupi_n_853,
     csa_tree_add_106_2_groupi_n_854, csa_tree_add_106_2_groupi_n_855,
     csa_tree_add_106_2_groupi_n_856, csa_tree_add_106_2_groupi_n_857,
     csa_tree_add_106_2_groupi_n_870, csa_tree_add_106_2_groupi_n_872,
     csa_tree_add_106_2_groupi_n_873, csa_tree_add_106_2_groupi_n_874,
     csa_tree_add_106_2_groupi_n_875, csa_tree_add_106_2_groupi_n_876,
     csa_tree_add_106_2_groupi_n_877, csa_tree_add_106_2_groupi_n_878,
     csa_tree_add_106_2_groupi_n_879, csa_tree_add_106_2_groupi_n_880,
     csa_tree_add_106_2_groupi_n_881, csa_tree_add_106_2_groupi_n_882,
     csa_tree_add_106_2_groupi_n_883, csa_tree_add_106_2_groupi_n_884,
     csa_tree_add_106_2_groupi_n_885, csa_tree_add_106_2_groupi_n_886,
     csa_tree_add_106_2_groupi_n_888, csa_tree_add_106_2_groupi_n_889,
     csa_tree_add_106_2_groupi_n_892, csa_tree_add_106_2_groupi_n_893,
     csa_tree_add_106_2_groupi_n_894, csa_tree_add_106_2_groupi_n_895,
     csa_tree_add_106_2_groupi_n_898, csa_tree_add_106_2_groupi_n_899,
     csa_tree_add_106_2_groupi_n_902, csa_tree_add_106_2_groupi_n_903,
     csa_tree_add_106_2_groupi_n_904, csa_tree_add_106_2_groupi_n_905,
     csa_tree_add_106_2_groupi_n_906, csa_tree_add_106_2_groupi_n_907,
     csa_tree_add_106_2_groupi_n_914, csa_tree_add_106_2_groupi_n_915,
     csa_tree_add_106_2_groupi_n_916, csa_tree_add_106_2_groupi_n_917,
     csa_tree_add_106_2_groupi_n_921, csa_tree_add_106_2_groupi_n_924,
     csa_tree_add_106_2_groupi_n_925, csa_tree_add_106_2_groupi_n_926,
     csa_tree_add_106_2_groupi_n_927, csa_tree_add_106_2_groupi_n_928,
     csa_tree_add_106_2_groupi_n_929, csa_tree_add_106_2_groupi_n_931,
     csa_tree_add_106_2_groupi_n_932, csa_tree_add_106_2_groupi_n_933,
     csa_tree_add_106_2_groupi_n_934, csa_tree_add_106_2_groupi_n_935,
     csa_tree_add_106_2_groupi_n_936, csa_tree_add_106_2_groupi_n_938,
     csa_tree_add_106_2_groupi_n_939, csa_tree_add_106_2_groupi_n_940,
     csa_tree_add_106_2_groupi_n_941, csa_tree_add_106_2_groupi_n_942,
     csa_tree_add_106_2_groupi_n_943, csa_tree_add_106_2_groupi_n_944,
     csa_tree_add_106_2_groupi_n_945, csa_tree_add_106_2_groupi_n_946,
     csa_tree_add_106_2_groupi_n_947, csa_tree_add_106_2_groupi_n_954,
     csa_tree_add_106_2_groupi_n_955, csa_tree_add_106_2_groupi_n_956,
     csa_tree_add_106_2_groupi_n_957, csa_tree_add_106_2_groupi_n_958,
     csa_tree_add_106_2_groupi_n_959, csa_tree_add_106_2_groupi_n_960,
     csa_tree_add_106_2_groupi_n_961, csa_tree_add_106_2_groupi_n_962,
     csa_tree_add_106_2_groupi_n_963, csa_tree_add_106_2_groupi_n_964,
     csa_tree_add_106_2_groupi_n_965, csa_tree_add_106_2_groupi_n_966,
     csa_tree_add_106_2_groupi_n_967, csa_tree_add_106_2_groupi_n_968,
     csa_tree_add_106_2_groupi_n_969, csa_tree_add_106_2_groupi_n_970,
     csa_tree_add_106_2_groupi_n_971, csa_tree_add_106_2_groupi_n_972,
     csa_tree_add_106_2_groupi_n_973, csa_tree_add_106_2_groupi_n_974,
     csa_tree_add_106_2_groupi_n_975, csa_tree_add_106_2_groupi_n_976,
     csa_tree_add_106_2_groupi_n_977, csa_tree_add_106_2_groupi_n_980,
     csa_tree_add_106_2_groupi_n_981, csa_tree_add_106_2_groupi_n_982,
     csa_tree_add_106_2_groupi_n_984, csa_tree_add_106_2_groupi_n_985,
     csa_tree_add_106_2_groupi_n_986, csa_tree_add_106_2_groupi_n_987,
     csa_tree_add_106_2_groupi_n_988, csa_tree_add_106_2_groupi_n_989,
     csa_tree_add_106_2_groupi_n_991, csa_tree_add_106_2_groupi_n_992,
     csa_tree_add_106_2_groupi_n_993, csa_tree_add_106_2_groupi_n_994,
     csa_tree_add_106_2_groupi_n_995, csa_tree_add_106_2_groupi_n_996,
     csa_tree_add_106_2_groupi_n_999, csa_tree_add_106_2_groupi_n_1000,
     csa_tree_add_106_2_groupi_n_1001, csa_tree_add_106_2_groupi_n_1002,
     csa_tree_add_106_2_groupi_n_1003, csa_tree_add_106_2_groupi_n_1004,
     csa_tree_add_106_2_groupi_n_1005, csa_tree_add_106_2_groupi_n_1006,
     csa_tree_add_106_2_groupi_n_1007, csa_tree_add_106_2_groupi_n_1008,
     csa_tree_add_106_2_groupi_n_1009, csa_tree_add_106_2_groupi_n_1010,
     csa_tree_add_106_2_groupi_n_1013, csa_tree_add_106_2_groupi_n_1014,
     csa_tree_add_106_2_groupi_n_1015, csa_tree_add_106_2_groupi_n_1016,
     csa_tree_add_106_2_groupi_n_1017, csa_tree_add_106_2_groupi_n_1018,
     csa_tree_add_106_2_groupi_n_1019, csa_tree_add_106_2_groupi_n_1020,
     csa_tree_add_106_2_groupi_n_1021, csa_tree_add_106_2_groupi_n_1022,
     csa_tree_add_106_2_groupi_n_1023, csa_tree_add_106_2_groupi_n_1024,
     csa_tree_add_106_2_groupi_n_1025, csa_tree_add_106_2_groupi_n_1027,
     csa_tree_add_106_2_groupi_n_1028, csa_tree_add_106_2_groupi_n_1029,
     csa_tree_add_106_2_groupi_n_1030, csa_tree_add_106_2_groupi_n_1031,
     csa_tree_add_106_2_groupi_n_1034, csa_tree_add_106_2_groupi_n_1035,
     csa_tree_add_106_2_groupi_n_1038, csa_tree_add_106_2_groupi_n_1039,
     csa_tree_add_106_2_groupi_n_1040, csa_tree_add_106_2_groupi_n_1041,
     csa_tree_add_106_2_groupi_n_1042, csa_tree_add_106_2_groupi_n_1043,
     csa_tree_add_106_2_groupi_n_1044, csa_tree_add_106_2_groupi_n_1047,
     csa_tree_add_106_2_groupi_n_1048, csa_tree_add_106_2_groupi_n_1049,
     csa_tree_add_106_2_groupi_n_1050, csa_tree_add_106_2_groupi_n_1051,
     csa_tree_add_106_2_groupi_n_1052, csa_tree_add_106_2_groupi_n_1053,
     csa_tree_add_106_2_groupi_n_1054, csa_tree_add_106_2_groupi_n_1057,
     csa_tree_add_106_2_groupi_n_1058, csa_tree_add_106_2_groupi_n_1063,
     csa_tree_add_106_2_groupi_n_1064, csa_tree_add_106_2_groupi_n_1067,
     csa_tree_add_106_2_groupi_n_1068, csa_tree_add_106_2_groupi_n_1069,
     csa_tree_add_106_2_groupi_n_1070, csa_tree_add_106_2_groupi_n_1071,
     csa_tree_add_106_2_groupi_n_1072, csa_tree_add_106_2_groupi_n_1073,
     csa_tree_add_106_2_groupi_n_1075, csa_tree_add_106_2_groupi_n_1076,
     csa_tree_add_106_2_groupi_n_1077, csa_tree_add_106_2_groupi_n_1078,
     csa_tree_add_106_2_groupi_n_1079, csa_tree_add_106_2_groupi_n_1080,
     csa_tree_add_106_2_groupi_n_1081, csa_tree_add_106_2_groupi_n_1082,
     csa_tree_add_106_2_groupi_n_1083, csa_tree_add_106_2_groupi_n_1084,
     csa_tree_add_106_2_groupi_n_1085, csa_tree_add_106_2_groupi_n_1086,
     csa_tree_add_106_2_groupi_n_1087, csa_tree_add_106_2_groupi_n_1088,
     csa_tree_add_106_2_groupi_n_1089, csa_tree_add_106_2_groupi_n_1090,
     csa_tree_add_106_2_groupi_n_1091, csa_tree_add_106_2_groupi_n_1094,
     csa_tree_add_106_2_groupi_n_1095, csa_tree_add_106_2_groupi_n_1096,
     csa_tree_add_106_2_groupi_n_1097, csa_tree_add_106_2_groupi_n_1098,
     csa_tree_add_106_2_groupi_n_1099, csa_tree_add_106_2_groupi_n_1100,
     csa_tree_add_106_2_groupi_n_1101, csa_tree_add_106_2_groupi_n_1102,
     csa_tree_add_106_2_groupi_n_1103, csa_tree_add_106_2_groupi_n_1106,
     csa_tree_add_106_2_groupi_n_1107, csa_tree_add_106_2_groupi_n_1108,
     csa_tree_add_106_2_groupi_n_1109, csa_tree_add_106_2_groupi_n_1110,
     csa_tree_add_106_2_groupi_n_1111, csa_tree_add_106_2_groupi_n_1112,
     csa_tree_add_106_2_groupi_n_1113, csa_tree_add_106_2_groupi_n_1114,
     csa_tree_add_106_2_groupi_n_1115, csa_tree_add_106_2_groupi_n_1118,
     csa_tree_add_106_2_groupi_n_1119, csa_tree_add_106_2_groupi_n_1120,
     csa_tree_add_106_2_groupi_n_1121, csa_tree_add_106_2_groupi_n_1150,
     csa_tree_add_106_2_groupi_n_1152, csa_tree_add_106_2_groupi_n_1154,
     csa_tree_add_106_2_groupi_n_1156, csa_tree_add_106_2_groupi_n_1158,
     csa_tree_add_106_2_groupi_n_1160, csa_tree_add_106_2_groupi_n_1162,
     csa_tree_mul_77_11_groupi_n_0, csa_tree_mul_77_11_groupi_n_1,
     csa_tree_mul_77_11_groupi_n_2, csa_tree_mul_77_11_groupi_n_3,
     csa_tree_mul_77_11_groupi_n_5, csa_tree_mul_77_11_groupi_n_6,
     csa_tree_mul_77_11_groupi_n_7, csa_tree_mul_77_11_groupi_n_9,
     csa_tree_mul_77_11_groupi_n_11, csa_tree_mul_77_11_groupi_n_12,
     csa_tree_mul_77_11_groupi_n_13, csa_tree_mul_77_11_groupi_n_14,
     csa_tree_mul_77_11_groupi_n_15, csa_tree_mul_77_11_groupi_n_16,
     csa_tree_mul_77_11_groupi_n_17, csa_tree_mul_77_11_groupi_n_18,
     csa_tree_mul_77_11_groupi_n_19, csa_tree_mul_77_11_groupi_n_20,
     csa_tree_mul_77_11_groupi_n_21, csa_tree_mul_77_11_groupi_n_22,
     csa_tree_mul_77_11_groupi_n_23, csa_tree_mul_77_11_groupi_n_24,
     csa_tree_mul_77_11_groupi_n_25, csa_tree_mul_77_11_groupi_n_26,
     csa_tree_mul_77_11_groupi_n_27, csa_tree_mul_77_11_groupi_n_28,
     csa_tree_mul_77_11_groupi_n_29, csa_tree_mul_77_11_groupi_n_30,
     csa_tree_mul_77_11_groupi_n_31, csa_tree_mul_77_11_groupi_n_32,
     csa_tree_mul_77_11_groupi_n_33, csa_tree_mul_77_11_groupi_n_34,
     csa_tree_mul_77_11_groupi_n_35, csa_tree_mul_77_11_groupi_n_36,
     csa_tree_mul_77_11_groupi_n_37, csa_tree_mul_77_11_groupi_n_38,
     csa_tree_mul_77_11_groupi_n_39, csa_tree_mul_77_11_groupi_n_40,
     csa_tree_mul_77_11_groupi_n_46, csa_tree_mul_77_11_groupi_n_47,
     csa_tree_mul_77_11_groupi_n_49, csa_tree_mul_77_11_groupi_n_50,
     csa_tree_mul_77_11_groupi_n_51, csa_tree_mul_77_11_groupi_n_52,
     csa_tree_mul_77_11_groupi_n_54, csa_tree_mul_77_11_groupi_n_55,
     csa_tree_mul_77_11_groupi_n_56, csa_tree_mul_77_11_groupi_n_57,
     csa_tree_mul_77_11_groupi_n_58, csa_tree_mul_77_11_groupi_n_59,
     csa_tree_mul_77_11_groupi_n_60, csa_tree_mul_77_11_groupi_n_61,
     csa_tree_mul_77_11_groupi_n_62, csa_tree_mul_77_11_groupi_n_63,
     csa_tree_mul_77_11_groupi_n_64, csa_tree_mul_77_11_groupi_n_65,
     csa_tree_mul_77_11_groupi_n_66, csa_tree_mul_77_11_groupi_n_67,
     csa_tree_mul_77_11_groupi_n_68, csa_tree_mul_77_11_groupi_n_69,
     csa_tree_mul_77_11_groupi_n_70, csa_tree_mul_77_11_groupi_n_71,
     csa_tree_mul_77_11_groupi_n_72, csa_tree_mul_77_11_groupi_n_73,
     csa_tree_mul_77_11_groupi_n_74, csa_tree_mul_77_11_groupi_n_75,
     csa_tree_mul_77_11_groupi_n_76, csa_tree_mul_77_11_groupi_n_77,
     csa_tree_mul_77_11_groupi_n_78, csa_tree_mul_77_11_groupi_n_79,
     csa_tree_mul_77_11_groupi_n_80, csa_tree_mul_77_11_groupi_n_81,
     csa_tree_mul_77_11_groupi_n_82, csa_tree_mul_77_11_groupi_n_83,
     csa_tree_mul_77_11_groupi_n_84, csa_tree_mul_77_11_groupi_n_85,
     csa_tree_mul_77_11_groupi_n_86, csa_tree_mul_77_11_groupi_n_87,
     csa_tree_mul_77_11_groupi_n_88, csa_tree_mul_77_11_groupi_n_89,
     csa_tree_mul_77_11_groupi_n_90, csa_tree_mul_77_11_groupi_n_91,
     csa_tree_mul_77_11_groupi_n_92, csa_tree_mul_77_11_groupi_n_93,
     csa_tree_mul_77_11_groupi_n_94, csa_tree_mul_77_11_groupi_n_95,
     csa_tree_mul_77_11_groupi_n_96, csa_tree_mul_77_11_groupi_n_97,
     csa_tree_mul_77_11_groupi_n_98, csa_tree_mul_77_11_groupi_n_99,
     csa_tree_mul_77_11_groupi_n_100, csa_tree_mul_77_11_groupi_n_101,
     csa_tree_mul_77_11_groupi_n_102, csa_tree_mul_77_11_groupi_n_103,
     csa_tree_mul_77_11_groupi_n_104, csa_tree_mul_77_11_groupi_n_105,
     csa_tree_mul_77_11_groupi_n_106, csa_tree_mul_77_11_groupi_n_107,
     csa_tree_mul_77_11_groupi_n_109, csa_tree_mul_77_11_groupi_n_110,
     csa_tree_mul_77_11_groupi_n_111, csa_tree_mul_77_11_groupi_n_112,
     csa_tree_mul_77_11_groupi_n_113, csa_tree_mul_77_11_groupi_n_114,
     csa_tree_mul_77_11_groupi_n_115, csa_tree_mul_77_11_groupi_n_116,
     csa_tree_mul_77_11_groupi_n_117, csa_tree_mul_77_11_groupi_n_118,
     csa_tree_mul_77_11_groupi_n_119, csa_tree_mul_77_11_groupi_n_120,
     csa_tree_mul_77_11_groupi_n_121, csa_tree_mul_77_11_groupi_n_122,
     csa_tree_mul_77_11_groupi_n_123, csa_tree_mul_77_11_groupi_n_124,
     csa_tree_mul_77_11_groupi_n_125, csa_tree_mul_77_11_groupi_n_126,
     csa_tree_mul_77_11_groupi_n_127, csa_tree_mul_77_11_groupi_n_128,
     csa_tree_mul_77_11_groupi_n_129, csa_tree_mul_77_11_groupi_n_130,
     csa_tree_mul_77_11_groupi_n_131, csa_tree_mul_77_11_groupi_n_132,
     csa_tree_mul_77_11_groupi_n_133, csa_tree_mul_77_11_groupi_n_134,
     csa_tree_mul_77_11_groupi_n_135, csa_tree_mul_77_11_groupi_n_136,
     csa_tree_mul_77_11_groupi_n_137, csa_tree_mul_77_11_groupi_n_138,
     csa_tree_mul_77_11_groupi_n_139, csa_tree_mul_77_11_groupi_n_140,
     csa_tree_mul_77_11_groupi_n_141, csa_tree_mul_77_11_groupi_n_142,
     csa_tree_mul_77_11_groupi_n_143, csa_tree_mul_77_11_groupi_n_144,
     csa_tree_mul_77_11_groupi_n_145, csa_tree_mul_77_11_groupi_n_146,
     csa_tree_mul_77_11_groupi_n_147, csa_tree_mul_77_11_groupi_n_148,
     csa_tree_mul_77_11_groupi_n_149, csa_tree_mul_77_11_groupi_n_150,
     csa_tree_mul_77_11_groupi_n_151, csa_tree_mul_77_11_groupi_n_152,
     csa_tree_mul_77_11_groupi_n_153, csa_tree_mul_77_11_groupi_n_154,
     csa_tree_mul_77_11_groupi_n_155, csa_tree_mul_77_11_groupi_n_156,
     csa_tree_mul_77_11_groupi_n_157, csa_tree_mul_77_11_groupi_n_158,
     csa_tree_mul_77_11_groupi_n_159, csa_tree_mul_77_11_groupi_n_160,
     csa_tree_mul_77_11_groupi_n_161, csa_tree_mul_77_11_groupi_n_162,
     csa_tree_mul_77_11_groupi_n_163, csa_tree_mul_77_11_groupi_n_164,
     csa_tree_mul_77_11_groupi_n_165, csa_tree_mul_77_11_groupi_n_166,
     csa_tree_mul_77_11_groupi_n_167, csa_tree_mul_77_11_groupi_n_168,
     csa_tree_mul_77_11_groupi_n_169, csa_tree_mul_77_11_groupi_n_170,
     csa_tree_mul_77_11_groupi_n_171, csa_tree_mul_77_11_groupi_n_172,
     csa_tree_mul_77_11_groupi_n_173, csa_tree_mul_77_11_groupi_n_174,
     csa_tree_mul_77_11_groupi_n_175, csa_tree_mul_77_11_groupi_n_176,
     csa_tree_mul_77_11_groupi_n_177, csa_tree_mul_77_11_groupi_n_178,
     csa_tree_mul_77_11_groupi_n_180, csa_tree_mul_77_11_groupi_n_181,
     csa_tree_mul_77_11_groupi_n_182, csa_tree_mul_77_11_groupi_n_183,
     csa_tree_mul_77_11_groupi_n_184, csa_tree_mul_77_11_groupi_n_185,
     csa_tree_mul_77_11_groupi_n_186, csa_tree_mul_77_11_groupi_n_187,
     csa_tree_mul_77_11_groupi_n_188, csa_tree_mul_77_11_groupi_n_189,
     csa_tree_mul_77_11_groupi_n_190, csa_tree_mul_77_11_groupi_n_191,
     csa_tree_mul_77_11_groupi_n_192, csa_tree_mul_77_11_groupi_n_193,
     csa_tree_mul_77_11_groupi_n_194, csa_tree_mul_77_11_groupi_n_195,
     csa_tree_mul_77_11_groupi_n_196, csa_tree_mul_77_11_groupi_n_197,
     csa_tree_mul_77_11_groupi_n_198, csa_tree_mul_77_11_groupi_n_199,
     csa_tree_mul_77_11_groupi_n_200, csa_tree_mul_77_11_groupi_n_201,
     csa_tree_mul_77_11_groupi_n_202, csa_tree_mul_77_11_groupi_n_203,
     csa_tree_mul_77_11_groupi_n_204, csa_tree_mul_77_11_groupi_n_205,
     csa_tree_mul_77_11_groupi_n_206, csa_tree_mul_77_11_groupi_n_207,
     csa_tree_mul_77_11_groupi_n_208, csa_tree_mul_77_11_groupi_n_209,
     csa_tree_mul_77_11_groupi_n_210, csa_tree_mul_77_11_groupi_n_211,
     csa_tree_mul_77_11_groupi_n_212, csa_tree_mul_77_11_groupi_n_213,
     csa_tree_mul_77_11_groupi_n_214, csa_tree_mul_77_11_groupi_n_215,
     csa_tree_mul_77_11_groupi_n_216, csa_tree_mul_77_11_groupi_n_217,
     csa_tree_mul_77_11_groupi_n_218, csa_tree_mul_77_11_groupi_n_219,
     csa_tree_mul_77_11_groupi_n_220, csa_tree_mul_77_11_groupi_n_221,
     csa_tree_mul_77_11_groupi_n_222, csa_tree_mul_77_11_groupi_n_223,
     csa_tree_mul_77_11_groupi_n_224, csa_tree_mul_77_11_groupi_n_225,
     csa_tree_mul_77_11_groupi_n_226, csa_tree_mul_77_11_groupi_n_227,
     csa_tree_mul_77_11_groupi_n_228, csa_tree_mul_77_11_groupi_n_229,
     csa_tree_mul_77_11_groupi_n_230, csa_tree_mul_77_11_groupi_n_231,
     csa_tree_mul_77_11_groupi_n_232, csa_tree_mul_77_11_groupi_n_233,
     csa_tree_mul_77_11_groupi_n_234, csa_tree_mul_77_11_groupi_n_235,
     csa_tree_mul_77_11_groupi_n_236, csa_tree_mul_77_11_groupi_n_237,
     csa_tree_mul_77_11_groupi_n_238, csa_tree_mul_77_11_groupi_n_239,
     csa_tree_mul_77_11_groupi_n_240, csa_tree_mul_77_11_groupi_n_241,
     csa_tree_mul_77_11_groupi_n_242, csa_tree_mul_77_11_groupi_n_243,
     csa_tree_mul_77_11_groupi_n_244, csa_tree_mul_77_11_groupi_n_245,
     csa_tree_mul_77_11_groupi_n_246, csa_tree_mul_77_11_groupi_n_247,
     csa_tree_mul_77_11_groupi_n_248, csa_tree_mul_77_11_groupi_n_249,
     csa_tree_mul_77_11_groupi_n_250, csa_tree_mul_77_11_groupi_n_251,
     csa_tree_mul_77_11_groupi_n_252, csa_tree_mul_77_11_groupi_n_253,
     csa_tree_mul_77_11_groupi_n_254, csa_tree_mul_77_11_groupi_n_255,
     csa_tree_mul_77_11_groupi_n_256, csa_tree_mul_77_11_groupi_n_257,
     csa_tree_mul_77_11_groupi_n_258, csa_tree_mul_77_11_groupi_n_259,
     csa_tree_mul_77_11_groupi_n_260, csa_tree_mul_77_11_groupi_n_261,
     csa_tree_mul_77_11_groupi_n_262, csa_tree_mul_77_11_groupi_n_263,
     csa_tree_mul_77_11_groupi_n_264, csa_tree_mul_77_11_groupi_n_265,
     csa_tree_mul_77_11_groupi_n_266, csa_tree_mul_77_11_groupi_n_267,
     csa_tree_mul_77_11_groupi_n_268, csa_tree_mul_77_11_groupi_n_269,
     csa_tree_mul_77_11_groupi_n_270, csa_tree_mul_77_11_groupi_n_271,
     csa_tree_mul_77_11_groupi_n_272, csa_tree_mul_77_11_groupi_n_273,
     csa_tree_mul_77_11_groupi_n_274, csa_tree_mul_77_11_groupi_n_275,
     csa_tree_mul_77_11_groupi_n_276, csa_tree_mul_77_11_groupi_n_277,
     csa_tree_mul_77_11_groupi_n_278, csa_tree_mul_77_11_groupi_n_279,
     csa_tree_mul_77_11_groupi_n_280, csa_tree_mul_77_11_groupi_n_281,
     csa_tree_mul_77_11_groupi_n_282, csa_tree_mul_77_11_groupi_n_283,
     csa_tree_mul_77_11_groupi_n_284, csa_tree_mul_77_11_groupi_n_285,
     csa_tree_mul_77_11_groupi_n_286, csa_tree_mul_77_11_groupi_n_287,
     csa_tree_mul_77_11_groupi_n_288, csa_tree_mul_77_11_groupi_n_289,
     csa_tree_mul_77_11_groupi_n_290, csa_tree_mul_77_11_groupi_n_291,
     csa_tree_mul_77_11_groupi_n_292, csa_tree_mul_77_11_groupi_n_293,
     csa_tree_mul_77_11_groupi_n_294, csa_tree_mul_77_11_groupi_n_295,
     csa_tree_mul_77_11_groupi_n_296, csa_tree_mul_77_11_groupi_n_297,
     csa_tree_mul_77_11_groupi_n_298, csa_tree_mul_77_11_groupi_n_299,
     csa_tree_mul_77_11_groupi_n_300, csa_tree_mul_77_11_groupi_n_301,
     csa_tree_mul_77_11_groupi_n_302, csa_tree_mul_77_11_groupi_n_303,
     csa_tree_mul_77_11_groupi_n_304, csa_tree_mul_77_11_groupi_n_305,
     csa_tree_mul_77_11_groupi_n_306, csa_tree_mul_77_11_groupi_n_307,
     csa_tree_mul_77_11_groupi_n_308, csa_tree_mul_77_11_groupi_n_309,
     csa_tree_mul_77_11_groupi_n_310, csa_tree_mul_77_11_groupi_n_311,
     csa_tree_mul_77_11_groupi_n_312, csa_tree_mul_77_11_groupi_n_313,
     csa_tree_mul_77_11_groupi_n_314, csa_tree_mul_77_11_groupi_n_316,
     csa_tree_mul_77_11_groupi_n_317, csa_tree_mul_77_11_groupi_n_318,
     csa_tree_mul_77_11_groupi_n_319, csa_tree_mul_77_11_groupi_n_320,
     csa_tree_mul_77_11_groupi_n_321, csa_tree_mul_77_11_groupi_n_322,
     csa_tree_mul_77_11_groupi_n_323, csa_tree_mul_77_11_groupi_n_324,
     csa_tree_mul_77_11_groupi_n_325, csa_tree_mul_77_11_groupi_n_326,
     csa_tree_mul_77_11_groupi_n_327, csa_tree_mul_77_11_groupi_n_328,
     csa_tree_mul_77_11_groupi_n_329, csa_tree_mul_77_11_groupi_n_330,
     csa_tree_mul_77_11_groupi_n_331, csa_tree_mul_77_11_groupi_n_332,
     csa_tree_mul_77_11_groupi_n_333, csa_tree_mul_77_11_groupi_n_334,
     csa_tree_mul_77_11_groupi_n_335, csa_tree_mul_77_11_groupi_n_338,
     csa_tree_mul_77_11_groupi_n_339, csa_tree_mul_77_11_groupi_n_342,
     csa_tree_mul_77_11_groupi_n_343, csa_tree_mul_77_11_groupi_n_344,
     csa_tree_mul_77_11_groupi_n_345, csa_tree_mul_77_11_groupi_n_346,
     csa_tree_mul_77_11_groupi_n_347, csa_tree_mul_77_11_groupi_n_349,
     csa_tree_mul_77_11_groupi_n_350, csa_tree_mul_77_11_groupi_n_351,
     csa_tree_mul_77_11_groupi_n_352, csa_tree_mul_77_11_groupi_n_353,
     csa_tree_mul_77_11_groupi_n_354, csa_tree_mul_77_11_groupi_n_355,
     csa_tree_mul_77_11_groupi_n_356, csa_tree_mul_77_11_groupi_n_357,
     csa_tree_mul_77_11_groupi_n_358, csa_tree_mul_77_11_groupi_n_359,
     csa_tree_mul_77_11_groupi_n_360, csa_tree_mul_77_11_groupi_n_361,
     csa_tree_mul_77_11_groupi_n_362, csa_tree_mul_77_11_groupi_n_363,
     csa_tree_mul_77_11_groupi_n_364, csa_tree_mul_77_11_groupi_n_365,
     csa_tree_mul_77_11_groupi_n_367, csa_tree_mul_77_11_groupi_n_368,
     csa_tree_mul_77_11_groupi_n_369, csa_tree_mul_77_11_groupi_n_371,
     csa_tree_mul_77_11_groupi_n_372, csa_tree_mul_77_11_groupi_n_373,
     csa_tree_mul_77_11_groupi_n_374, csa_tree_mul_77_11_groupi_n_377,
     csa_tree_mul_77_11_groupi_n_378, csa_tree_mul_77_11_groupi_n_379,
     csa_tree_mul_77_11_groupi_n_380, csa_tree_mul_77_11_groupi_n_381,
     csa_tree_mul_77_11_groupi_n_383, csa_tree_mul_77_11_groupi_n_384,
     csa_tree_mul_77_11_groupi_n_385, csa_tree_mul_77_11_groupi_n_386,
     csa_tree_mul_77_11_groupi_n_387, csa_tree_mul_77_11_groupi_n_388,
     csa_tree_mul_77_11_groupi_n_389, csa_tree_mul_77_11_groupi_n_395,
     csa_tree_mul_77_11_groupi_n_396, csa_tree_mul_77_11_groupi_n_397,
     csa_tree_mul_77_11_groupi_n_398, csa_tree_mul_77_11_groupi_n_401,
     csa_tree_mul_77_11_groupi_n_402, csa_tree_mul_77_11_groupi_n_403,
     csa_tree_mul_77_11_groupi_n_404, csa_tree_mul_77_11_groupi_n_405,
     csa_tree_mul_77_11_groupi_n_406, csa_tree_mul_77_11_groupi_n_407,
     csa_tree_mul_77_11_groupi_n_408, csa_tree_mul_77_11_groupi_n_409,
     csa_tree_mul_77_11_groupi_n_412, csa_tree_mul_77_11_groupi_n_413,
     csa_tree_mul_77_11_groupi_n_414, csa_tree_mul_77_11_groupi_n_416,
     csa_tree_mul_77_11_groupi_n_417, csa_tree_mul_77_11_groupi_n_418,
     csa_tree_mul_77_11_groupi_n_419, csa_tree_mul_77_11_groupi_n_420,
     csa_tree_mul_77_11_groupi_n_421, csa_tree_mul_77_11_groupi_n_422,
     csa_tree_mul_77_11_groupi_n_423, csa_tree_mul_77_11_groupi_n_424,
     csa_tree_mul_77_11_groupi_n_425, csa_tree_mul_77_11_groupi_n_426,
     csa_tree_mul_77_11_groupi_n_427, csa_tree_mul_77_11_groupi_n_428,
     csa_tree_mul_77_11_groupi_n_429, csa_tree_mul_77_11_groupi_n_430,
     csa_tree_mul_77_11_groupi_n_433, csa_tree_mul_77_11_groupi_n_434,
     csa_tree_mul_77_11_groupi_n_435, csa_tree_mul_77_11_groupi_n_438,
     csa_tree_mul_77_11_groupi_n_439, csa_tree_mul_77_11_groupi_n_440,
     csa_tree_mul_77_11_groupi_n_441, csa_tree_mul_77_11_groupi_n_442,
     csa_tree_mul_77_11_groupi_n_444, csa_tree_mul_77_11_groupi_n_445,
     csa_tree_mul_77_11_groupi_n_447, csa_tree_mul_77_11_groupi_n_448,
     csa_tree_mul_77_11_groupi_n_449, csa_tree_mul_77_11_groupi_n_450,
     csa_tree_mul_77_11_groupi_n_451, csa_tree_mul_77_11_groupi_n_452,
     csa_tree_mul_77_11_groupi_n_453, csa_tree_mul_77_11_groupi_n_454,
     csa_tree_mul_77_11_groupi_n_455, csa_tree_mul_77_11_groupi_n_457,
     csa_tree_mul_77_11_groupi_n_459, csa_tree_mul_77_11_groupi_n_460,
     csa_tree_mul_77_11_groupi_n_461, csa_tree_mul_77_11_groupi_n_462,
     csa_tree_mul_77_11_groupi_n_463, csa_tree_mul_77_11_groupi_n_464,
     csa_tree_mul_77_11_groupi_n_469, csa_tree_mul_77_11_groupi_n_471,
     csa_tree_mul_77_11_groupi_n_472, csa_tree_mul_77_11_groupi_n_473,
     csa_tree_mul_77_11_groupi_n_474, csa_tree_mul_77_11_groupi_n_475,
     csa_tree_mul_77_11_groupi_n_476, csa_tree_mul_77_11_groupi_n_477,
     csa_tree_mul_77_11_groupi_n_478, csa_tree_mul_77_11_groupi_n_479,
     csa_tree_mul_77_11_groupi_n_480, csa_tree_mul_77_11_groupi_n_481,
     csa_tree_mul_77_11_groupi_n_483, csa_tree_mul_77_11_groupi_n_484,
     csa_tree_mul_77_11_groupi_n_485, csa_tree_mul_77_11_groupi_n_486,
     csa_tree_mul_77_11_groupi_n_487, csa_tree_mul_77_11_groupi_n_488,
     csa_tree_mul_77_11_groupi_n_489, csa_tree_mul_77_11_groupi_n_490,
     csa_tree_mul_77_11_groupi_n_492, csa_tree_mul_77_11_groupi_n_493,
     csa_tree_mul_77_11_groupi_n_494, csa_tree_mul_77_11_groupi_n_495,
     csa_tree_mul_77_11_groupi_n_497, csa_tree_mul_77_11_groupi_n_498,
     csa_tree_mul_77_11_groupi_n_499, csa_tree_mul_77_11_groupi_n_500,
     csa_tree_mul_77_11_groupi_n_501, csa_tree_mul_77_11_groupi_n_503,
     csa_tree_mul_77_11_groupi_n_504, csa_tree_mul_77_11_groupi_n_505,
     csa_tree_mul_77_11_groupi_n_506, csa_tree_mul_77_11_groupi_n_507,
     csa_tree_mul_77_11_groupi_n_508, csa_tree_mul_77_11_groupi_n_509,
     csa_tree_mul_77_11_groupi_n_510, csa_tree_mul_77_11_groupi_n_511,
     csa_tree_mul_77_11_groupi_n_512, csa_tree_mul_77_11_groupi_n_513,
     csa_tree_mul_77_11_groupi_n_514, csa_tree_mul_77_11_groupi_n_515,
     csa_tree_mul_77_11_groupi_n_517, csa_tree_mul_77_11_groupi_n_518,
     csa_tree_mul_77_11_groupi_n_520, csa_tree_mul_77_11_groupi_n_521,
     csa_tree_mul_77_11_groupi_n_522, csa_tree_mul_77_11_groupi_n_523,
     csa_tree_mul_77_11_groupi_n_524, csa_tree_mul_77_11_groupi_n_525,
     csa_tree_mul_77_11_groupi_n_526, csa_tree_mul_77_11_groupi_n_527,
     csa_tree_mul_77_11_groupi_n_528, csa_tree_mul_77_11_groupi_n_530,
     csa_tree_mul_77_11_groupi_n_531, csa_tree_mul_77_11_groupi_n_533,
     csa_tree_mul_77_11_groupi_n_534, csa_tree_mul_77_11_groupi_n_535,
     csa_tree_mul_77_11_groupi_n_536, csa_tree_mul_77_11_groupi_n_537,
     csa_tree_mul_77_11_groupi_n_538, csa_tree_mul_77_11_groupi_n_539,
     csa_tree_mul_77_11_groupi_n_542, csa_tree_mul_77_11_groupi_n_544,
     csa_tree_mul_77_11_groupi_n_545, csa_tree_mul_77_11_groupi_n_546,
     csa_tree_mul_77_11_groupi_n_547, csa_tree_mul_77_11_groupi_n_548,
     csa_tree_mul_77_11_groupi_n_549, csa_tree_mul_77_11_groupi_n_550,
     csa_tree_mul_77_11_groupi_n_551, csa_tree_mul_77_11_groupi_n_552,
     csa_tree_mul_77_11_groupi_n_553, csa_tree_mul_77_11_groupi_n_554,
     csa_tree_mul_77_11_groupi_n_555, csa_tree_mul_77_11_groupi_n_556,
     csa_tree_mul_77_11_groupi_n_557, csa_tree_mul_77_11_groupi_n_559,
     csa_tree_mul_77_11_groupi_n_560, csa_tree_mul_77_11_groupi_n_561,
     csa_tree_mul_77_11_groupi_n_563, csa_tree_mul_77_11_groupi_n_564,
     csa_tree_mul_77_11_groupi_n_565, csa_tree_mul_77_11_groupi_n_566,
     csa_tree_mul_77_11_groupi_n_567, csa_tree_mul_77_11_groupi_n_568,
     csa_tree_mul_77_11_groupi_n_570, csa_tree_mul_77_11_groupi_n_571,
     csa_tree_mul_77_11_groupi_n_572, csa_tree_mul_77_11_groupi_n_573,
     csa_tree_mul_77_11_groupi_n_574, csa_tree_mul_77_11_groupi_n_575,
     csa_tree_mul_77_11_groupi_n_576, csa_tree_mul_77_11_groupi_n_581,
     csa_tree_mul_77_11_groupi_n_582, csa_tree_mul_77_11_groupi_n_583,
     csa_tree_mul_77_11_groupi_n_584, csa_tree_mul_77_11_groupi_n_585,
     csa_tree_mul_77_11_groupi_n_586, csa_tree_mul_77_11_groupi_n_587,
     csa_tree_mul_77_11_groupi_n_590, csa_tree_mul_77_11_groupi_n_591,
     csa_tree_mul_77_11_groupi_n_592, csa_tree_mul_77_11_groupi_n_593,
     csa_tree_mul_77_11_groupi_n_594, csa_tree_mul_77_11_groupi_n_600,
     csa_tree_mul_77_11_groupi_n_601, csa_tree_mul_77_11_groupi_n_603,
     csa_tree_mul_77_11_groupi_n_604, csa_tree_mul_77_11_groupi_n_605,
     csa_tree_mul_77_11_groupi_n_606, csa_tree_mul_77_11_groupi_n_607,
     csa_tree_mul_77_11_groupi_n_608, csa_tree_mul_77_11_groupi_n_609,
     csa_tree_mul_77_11_groupi_n_613, csa_tree_mul_77_11_groupi_n_614,
     csa_tree_mul_77_11_groupi_n_615, csa_tree_mul_77_11_groupi_n_617,
     csa_tree_mul_77_11_groupi_n_619, csa_tree_mul_77_11_groupi_n_620,
     csa_tree_mul_77_11_groupi_n_621, final_adder_add_69_2_n_2,
     final_adder_add_69_2_n_4, final_adder_add_69_2_n_6,
     final_adder_add_69_2_n_8, final_adder_add_69_2_n_10,
     final_adder_add_69_2_n_12, final_adder_add_86_2_n_1,
     final_adder_add_86_2_n_3, final_adder_add_86_2_n_19,
     final_adder_add_86_2_n_21, final_adder_add_86_2_n_23,
     final_adder_add_86_2_n_25, final_adder_add_86_2_n_27,
     final_adder_add_86_2_n_29, final_adder_add_86_2_n_31,
     final_adder_add_86_2_n_33, final_adder_add_86_2_n_35,
     final_adder_add_86_2_n_37, final_adder_add_86_2_n_39,
     final_adder_add_86_2_n_41, final_adder_add_86_2_n_43,
     final_adder_add_86_2_n_45, final_adder_add_86_2_n_47,
     final_adder_add_86_2_n_49, mul_74_11_n_0, mul_74_11_n_2, mul_74_11_n_4,
     mul_74_11_n_5, mul_74_11_n_6, mul_74_11_n_7, mul_74_11_n_8, mul_74_11_n_9,
     mul_74_11_n_10, mul_74_11_n_11, mul_74_11_n_12, mul_74_11_n_13,
     mul_74_11_n_14, mul_74_11_n_15, mul_74_11_n_16, mul_74_11_n_17,
     mul_74_11_n_18, mul_74_11_n_19, mul_74_11_n_20, mul_74_11_n_21,
     mul_74_11_n_22, mul_74_11_n_23, mul_74_11_n_24, mul_74_11_n_25,
     mul_74_11_n_26, mul_74_11_n_27, mul_74_11_n_28, mul_74_11_n_29,
     mul_74_11_n_30, mul_74_11_n_31, mul_74_11_n_33, mul_74_11_n_34,
     mul_74_11_n_35, mul_74_11_n_36, mul_74_11_n_37, mul_74_11_n_38,
     mul_74_11_n_39, mul_74_11_n_40, mul_74_11_n_41, mul_74_11_n_42,
     mul_74_11_n_43, mul_74_11_n_44, mul_74_11_n_45, mul_74_11_n_46,
     mul_74_11_n_47, mul_74_11_n_48, mul_74_11_n_49, mul_74_11_n_50,
     mul_74_11_n_51, mul_74_11_n_52, mul_74_11_n_53, mul_74_11_n_68,
     mul_74_11_n_78, mul_74_11_n_84, mul_74_11_n_85, mul_74_11_n_86,
     mul_74_11_n_87, mul_74_11_n_88, mul_74_11_n_89, mul_74_11_n_90,
     mul_74_11_n_91, mul_74_11_n_92, mul_74_11_n_93, mul_74_11_n_94,
     mul_74_11_n_98, mul_74_11_n_99, mul_74_11_n_100, mul_74_11_n_101,
     mul_74_11_n_102, mul_74_11_n_108, mul_74_11_n_109, mul_74_11_n_110,
     mul_74_11_n_115, mul_74_11_n_117, mul_74_11_n_118, mul_74_11_n_119,
     mul_74_11_n_120, mul_74_11_n_121, mul_74_11_n_122, mul_74_11_n_123,
     mul_74_11_n_125, mul_74_11_n_126, mul_74_11_n_128, mul_74_11_n_130,
     mul_74_11_n_133, mul_74_11_n_134, mul_74_11_n_138, mul_74_11_n_139,
     mul_74_11_n_140, mul_74_11_n_141, mul_74_11_n_143, mul_74_11_n_146,
     mul_74_11_n_153, mul_74_11_n_154, mul_74_11_n_155, mul_74_11_n_156,
     mul_74_11_n_157, mul_74_11_n_159, mul_74_11_n_160, mul_74_11_n_162,
     mul_74_11_n_163, mul_74_11_n_164, mul_74_11_n_165, mul_74_11_n_166,
     mul_74_11_n_167, mul_74_11_n_169, mul_74_11_n_170, mul_74_11_n_171,
     mul_74_11_n_173, mul_74_11_n_174, mul_74_11_n_175, mul_74_11_n_176,
     mul_74_11_n_177, mul_74_11_n_178, mul_74_11_n_179, mul_74_11_n_180,
     mul_74_11_n_181, mul_74_11_n_184, mul_74_11_n_186, mul_74_11_n_189,
     mul_74_11_n_191, mul_74_11_n_192, mul_74_11_n_193, mul_74_11_n_194,
     mul_74_11_n_195, mul_74_11_n_196, mul_74_11_n_197, mul_74_11_n_198,
     mul_74_11_n_199, mul_74_11_n_200, mul_74_11_n_201, mul_74_11_n_202,
     mul_74_11_n_203, mul_74_11_n_204, mul_74_11_n_205, mul_74_11_n_206,
     mul_74_11_n_207, mul_74_11_n_208, mul_74_11_n_209, mul_74_11_n_210,
     mul_74_11_n_211, mul_74_11_n_212, mul_74_11_n_213, mul_74_11_n_215,
     mul_74_11_n_216, mul_74_11_n_217, mul_74_11_n_218, mul_74_11_n_219,
     mul_74_11_n_220, mul_74_11_n_221, mul_74_11_n_222, mul_74_11_n_223,
     mul_74_11_n_224, mul_74_11_n_225, mul_74_11_n_226, mul_74_11_n_227,
     mul_74_11_n_228, mul_74_11_n_229, mul_74_11_n_230, mul_74_11_n_231,
     mul_74_11_n_232, mul_74_11_n_233, mul_74_11_n_234, mul_74_11_n_235,
     mul_74_11_n_236, mul_74_11_n_237, mul_74_11_n_238, mul_74_11_n_239,
     mul_74_11_n_240, mul_74_11_n_241, mul_74_11_n_242, mul_74_11_n_243,
     mul_74_11_n_244, mul_74_11_n_245, mul_74_11_n_246, mul_74_11_n_247,
     mul_74_11_n_248, mul_74_11_n_249, mul_74_11_n_250, mul_74_11_n_251,
     mul_74_11_n_252, mul_74_11_n_253, mul_74_11_n_254, mul_74_11_n_255,
     mul_74_11_n_257, mul_74_11_n_258, mul_74_11_n_259, mul_74_11_n_260,
     mul_74_11_n_261, mul_74_11_n_262, mul_74_11_n_263, mul_74_11_n_264,
     mul_74_11_n_265, mul_74_11_n_266, mul_74_11_n_267, mul_74_11_n_268,
     mul_74_11_n_269, mul_74_11_n_270, mul_74_11_n_271, mul_74_11_n_272,
     mul_74_11_n_273, mul_74_11_n_274, mul_74_11_n_275, mul_74_11_n_276,
     mul_74_11_n_277, mul_74_11_n_278, mul_74_11_n_279, mul_74_11_n_280,
     mul_74_11_n_281, mul_74_11_n_282, mul_74_11_n_283, mul_74_11_n_284,
     mul_74_11_n_285, mul_74_11_n_286, mul_74_11_n_287, mul_74_11_n_288,
     mul_74_11_n_289, mul_74_11_n_290, mul_74_11_n_291, mul_74_11_n_292,
     mul_74_11_n_293, mul_74_11_n_294, mul_74_11_n_295, mul_74_11_n_296,
     mul_74_11_n_297, mul_74_11_n_298, mul_74_11_n_299, mul_74_11_n_300,
     mul_74_11_n_301, mul_74_11_n_302, mul_74_11_n_303, mul_74_11_n_304,
     mul_74_11_n_305, mul_74_11_n_306, mul_74_11_n_307, mul_74_11_n_308,
     mul_74_11_n_309, mul_74_11_n_310, mul_74_11_n_311, mul_74_11_n_312,
     mul_74_11_n_313, mul_74_11_n_314, mul_74_11_n_315, mul_74_11_n_316,
     mul_74_11_n_317, mul_74_11_n_318, mul_74_11_n_319, mul_74_11_n_320,
     mul_74_11_n_321, mul_74_11_n_322, mul_74_11_n_323, mul_74_11_n_324,
     mul_74_11_n_325, mul_74_11_n_326, mul_74_11_n_327, mul_74_11_n_328,
     mul_74_11_n_329, mul_74_11_n_330, mul_74_11_n_331, mul_74_11_n_332,
     mul_74_11_n_333, mul_74_11_n_334, mul_74_11_n_335, mul_74_11_n_336,
     mul_74_11_n_339, mul_74_11_n_340, mul_74_11_n_341, mul_74_11_n_342,
     mul_74_11_n_343, mul_74_11_n_344, mul_74_11_n_345, mul_74_11_n_346,
     mul_74_11_n_347, mul_74_11_n_348, mul_74_11_n_349, mul_74_11_n_350,
     mul_74_11_n_351, mul_74_11_n_352, mul_74_11_n_353, mul_74_11_n_354,
     mul_74_11_n_355, mul_74_11_n_356, mul_74_11_n_357, mul_74_11_n_360,
     mul_74_11_n_362, mul_74_11_n_364, mul_74_11_n_366, mul_74_11_n_367,
     mul_74_11_n_368, mul_74_11_n_369, mul_74_11_n_370, mul_74_11_n_371,
     mul_74_11_n_372, mul_74_11_n_373, mul_74_11_n_374, mul_74_11_n_375,
     mul_74_11_n_376, mul_74_11_n_377, mul_74_11_n_378, mul_74_11_n_379,
     mul_74_11_n_380, mul_74_11_n_381, mul_74_11_n_382, mul_74_11_n_383,
     mul_74_11_n_384, mul_74_11_n_385, mul_74_11_n_386, mul_74_11_n_387,
     mul_74_11_n_388, mul_74_11_n_389, mul_74_11_n_390, mul_74_11_n_391,
     mul_74_11_n_392, mul_74_11_n_393, mul_74_11_n_394, mul_74_11_n_395,
     mul_74_11_n_396, mul_74_11_n_397, mul_74_11_n_398, mul_74_11_n_399,
     mul_74_11_n_400, mul_74_11_n_401, mul_74_11_n_402, mul_74_11_n_403,
     mul_74_11_n_404, mul_74_11_n_405, mul_74_11_n_406, mul_74_11_n_407,
     mul_74_11_n_408, mul_74_11_n_409, mul_74_11_n_410, mul_74_11_n_412,
     mul_74_11_n_413, mul_74_11_n_414, mul_74_11_n_415, mul_74_11_n_416,
     mul_74_11_n_417, mul_74_11_n_418, mul_74_11_n_419, mul_74_11_n_420,
     mul_74_11_n_421, mul_74_11_n_422, mul_74_11_n_423, mul_74_11_n_424,
     mul_74_11_n_425, mul_74_11_n_426, mul_74_11_n_427, mul_74_11_n_428,
     mul_74_11_n_429, mul_74_11_n_430, mul_74_11_n_431, mul_74_11_n_432,
     mul_74_11_n_433, mul_74_11_n_434, mul_74_11_n_435, mul_74_11_n_436,
     mul_74_11_n_437, mul_74_11_n_438, mul_74_11_n_439, mul_74_11_n_440,
     mul_74_11_n_441, mul_74_11_n_442, mul_74_11_n_443, mul_74_11_n_444,
     mul_74_11_n_445, mul_74_11_n_446, mul_74_11_n_448, mul_74_11_n_449,
     mul_74_11_n_450, mul_74_11_n_451, mul_74_11_n_452, mul_74_11_n_453,
     mul_74_11_n_454, mul_74_11_n_455, mul_74_11_n_456, mul_74_11_n_457,
     mul_74_11_n_458, mul_74_11_n_459, mul_74_11_n_460, mul_74_11_n_461,
     mul_74_11_n_462, mul_74_11_n_464, mul_74_11_n_465, mul_74_11_n_468,
     mul_74_11_n_469, mul_74_11_n_470, mul_74_11_n_471, mul_74_11_n_472,
     mul_74_11_n_476, mul_74_11_n_477, mul_74_11_n_478, mul_74_11_n_479,
     mul_74_11_n_480, mul_74_11_n_481, mul_74_11_n_482, mul_74_11_n_483,
     mul_74_11_n_484, mul_74_11_n_485, mul_74_11_n_489, mul_74_11_n_490,
     mul_74_11_n_491, mul_74_11_n_492, mul_74_11_n_493, mul_74_11_n_495,
     mul_74_11_n_496, mul_74_11_n_497, mul_74_11_n_498, mul_74_11_n_499,
     mul_74_11_n_500, mul_74_11_n_501, mul_74_11_n_502, mul_74_11_n_503,
     mul_74_11_n_504, mul_74_11_n_505, mul_74_11_n_506, mul_74_11_n_507,
     mul_74_11_n_508, mul_74_11_n_509, mul_74_11_n_510, mul_74_11_n_512,
     mul_74_11_n_513, mul_74_11_n_516, mul_74_11_n_517, mul_74_11_n_518,
     mul_74_11_n_519, mul_74_11_n_520, mul_74_11_n_522, mul_74_11_n_523,
     mul_74_11_n_524, mul_74_11_n_525, mul_74_11_n_526, mul_74_11_n_527,
     mul_74_11_n_528, mul_74_11_n_529, mul_74_11_n_530, mul_74_11_n_531,
     mul_74_11_n_532, mul_74_11_n_533, mul_74_11_n_534, mul_74_11_n_535,
     mul_74_11_n_536, mul_74_11_n_537, mul_74_11_n_538, mul_74_11_n_539,
     mul_74_11_n_540, mul_74_11_n_542, mul_74_11_n_543, mul_74_11_n_545,
     mul_74_11_n_546, mul_74_11_n_547, mul_74_11_n_548, mul_74_11_n_549,
     mul_74_11_n_550, mul_74_11_n_551, mul_74_11_n_552, mul_74_11_n_554,
     mul_74_11_n_555, mul_74_11_n_556, mul_74_11_n_558, mul_74_11_n_559,
     mul_74_11_n_560, mul_74_11_n_561, mul_74_11_n_564, mul_74_11_n_566,
     mul_74_11_n_568, mul_74_11_n_570, mul_109_11_n_0, mul_109_11_n_1,
     mul_109_11_n_2, mul_109_11_n_3, mul_109_11_n_12, mul_109_11_n_13,
     mul_109_11_n_14, mul_109_11_n_15, mul_109_11_n_16, mul_109_11_n_17,
     mul_109_11_n_19, mul_109_11_n_25, mul_109_11_n_26, mul_109_11_n_28,
     mul_109_11_n_31, mul_109_11_n_38, mul_109_11_n_39, mul_109_11_n_41,
     mul_109_11_n_43, mul_109_11_n_52, mul_109_11_n_56, mul_109_11_n_61,
     mul_109_11_n_62, mul_109_11_n_63, mul_109_11_n_64, mul_109_11_n_65,
     mul_109_11_n_69, mul_109_11_n_72, mul_109_11_n_73, mul_109_11_n_74,
     mul_109_11_n_75, mul_109_11_n_76, mul_109_11_n_77, mul_109_11_n_78,
     mul_109_11_n_79, mul_109_11_n_81, mul_109_11_n_82, mul_109_11_n_83,
     mul_109_11_n_84, mul_109_11_n_85, mul_109_11_n_86, mul_109_11_n_87,
     mul_109_11_n_88, mul_109_11_n_89, mul_109_11_n_90, mul_109_11_n_92,
     mul_109_11_n_93, mul_109_11_n_94, mul_109_11_n_95, mul_109_11_n_96,
     mul_109_11_n_98, mul_109_11_n_99, mul_109_11_n_100, mul_109_11_n_101,
     mul_109_11_n_102, mul_109_11_n_103, mul_109_11_n_104, mul_109_11_n_105,
     mul_109_11_n_106, mul_109_11_n_107, mul_109_11_n_108, mul_109_11_n_109,
     mul_109_11_n_110, mul_109_11_n_111, mul_109_11_n_112, mul_109_11_n_113,
     mul_109_11_n_114, mul_109_11_n_115, mul_109_11_n_116, mul_109_11_n_117,
     mul_109_11_n_118, mul_109_11_n_119, mul_109_11_n_120, mul_109_11_n_121,
     mul_109_11_n_122, mul_109_11_n_123, mul_109_11_n_124, mul_109_11_n_125,
     mul_109_11_n_126, mul_109_11_n_127, mul_109_11_n_128, mul_109_11_n_129,
     mul_109_11_n_130, mul_109_11_n_131, mul_109_11_n_132, mul_109_11_n_133,
     mul_109_11_n_134, mul_109_11_n_135, mul_109_11_n_136, mul_109_11_n_137,
     mul_109_11_n_138, mul_109_11_n_139, mul_109_11_n_140, mul_109_11_n_142,
     mul_109_11_n_143, mul_109_11_n_144, mul_109_11_n_145, mul_109_11_n_146,
     mul_109_11_n_147, mul_109_11_n_148, mul_109_11_n_149, mul_109_11_n_151,
     mul_109_11_n_153, mul_109_11_n_154, mul_109_11_n_157, mul_109_11_n_158,
     mul_109_11_n_159, mul_109_11_n_161, mul_109_11_n_162, mul_109_11_n_163,
     mul_109_11_n_164, mul_109_11_n_165, mul_109_11_n_167, mul_109_11_n_168,
     mul_109_11_n_169, mul_109_11_n_170, mul_109_11_n_171, mul_109_11_n_172,
     mul_109_11_n_173, mul_109_11_n_174, mul_109_11_n_177, mul_109_11_n_178,
     mul_109_11_n_183, mul_109_11_n_184, mul_109_11_n_187, mul_109_11_n_188,
     mul_109_11_n_189, mul_109_11_n_190, mul_109_11_n_191, mul_109_11_n_192,
     mul_109_11_n_193, mul_109_11_n_194, mul_109_11_n_195, mul_109_11_n_196,
     mul_109_11_n_199, mul_109_11_n_200, mul_109_11_n_206, mul_109_11_n_207,
     mul_109_11_n_208, mul_109_11_n_209, mul_109_11_n_210, mul_109_11_n_211,
     mul_109_11_n_212, mul_109_11_n_213, mul_109_11_n_214, mul_109_11_n_215,
     mul_109_11_n_221, mul_109_11_n_223, mul_109_11_n_224, mul_109_11_n_225,
     mul_109_11_n_226, mul_109_11_n_227, mul_109_11_n_228, mul_109_11_n_230,
     mul_109_11_n_231, mul_109_11_n_232, mul_109_11_n_233, mul_109_11_n_234,
     mul_109_11_n_235, mul_109_11_n_236, mul_109_11_n_237, mul_109_11_n_238,
     mul_109_11_n_239, mul_109_11_n_240, mul_109_11_n_241, mul_109_11_n_242,
     mul_109_11_n_245, mul_109_11_n_246, mul_109_11_n_247, mul_109_11_n_250,
     mul_109_11_n_252, mul_109_11_n_255, mul_109_11_n_256, mul_109_11_n_257,
     mul_109_11_n_258, mul_109_11_n_259, mul_109_11_n_260, mul_109_11_n_261,
     mul_109_11_n_262, mul_109_11_n_263, mul_109_11_n_264, mul_109_11_n_265,
     mul_109_11_n_266, mul_109_11_n_267, mul_109_11_n_268, mul_109_11_n_271,
     mul_109_11_n_272, mul_109_11_n_275, mul_109_11_n_276, mul_109_11_n_277,
     mul_109_11_n_278, mul_109_11_n_279, mul_109_11_n_280, mul_109_11_n_281,
     mul_109_11_n_282, mul_109_11_n_285, mul_109_11_n_286, mul_109_11_n_287,
     mul_109_11_n_288, mul_109_11_n_294, mul_109_11_n_295, mul_109_11_n_296,
     mul_109_11_n_297, mul_109_11_n_298, mul_109_11_n_301, mul_109_11_n_302,
     mul_109_11_n_303, mul_109_11_n_304, mul_109_11_n_305, mul_109_11_n_306,
     mul_109_11_n_307, mul_109_11_n_312, mul_109_11_n_313, mul_109_11_n_316,
     mul_109_11_n_317, mul_109_11_n_318, mul_109_11_n_320, mul_109_11_n_321,
     mul_109_11_n_322, mul_109_11_n_327, mul_109_11_n_328, mul_109_11_n_329,
     mul_109_11_n_332, mul_109_11_n_333, mul_109_11_n_334, mul_109_11_n_335,
     mul_109_11_n_340, mul_109_11_n_341, mul_109_11_n_344, mul_109_11_n_345,
     mul_109_11_n_346, mul_109_11_n_347, mul_109_11_n_348, mul_109_11_n_352,
     mul_109_11_n_353, mul_109_11_n_356, mul_109_11_n_357, mul_109_11_n_360,
     mul_109_11_n_361, mul_109_11_n_364, mul_109_11_n_365, mul_109_11_n_366,
     mul_109_11_n_367, mul_109_11_n_370, mul_109_11_n_371, mul_109_11_n_372,
     mul_109_11_n_374, mul_109_11_n_375, mul_109_11_n_376, mul_109_11_n_377,
     mul_109_11_n_378, mul_109_11_n_379, mul_109_11_n_380, mul_109_11_n_381,
     mul_109_11_n_382, mul_109_11_n_383, mul_109_11_n_384, mul_109_11_n_385,
     mul_109_11_n_386, mul_109_11_n_387, mul_109_11_n_388, mul_109_11_n_389,
     mul_109_11_n_390, mul_109_11_n_391, mul_109_11_n_392, mul_109_11_n_393,
     mul_109_11_n_394, mul_109_11_n_395, mul_109_11_n_396, mul_109_11_n_397,
     mul_109_11_n_398, mul_109_11_n_399, mul_109_11_n_400, mul_109_11_n_401,
     mul_109_11_n_402, mul_109_11_n_403, mul_109_11_n_404, mul_109_11_n_405,
     mul_109_11_n_406, mul_109_11_n_407, mul_109_11_n_408, mul_109_11_n_409,
     mul_109_11_n_410, mul_109_11_n_411, mul_109_11_n_412, mul_109_11_n_413,
     mul_109_11_n_414, mul_109_11_n_415, mul_109_11_n_416, mul_109_11_n_417,
     mul_109_11_n_418, mul_109_11_n_419, mul_109_11_n_420, mul_109_11_n_421,
     mul_109_11_n_422, mul_109_11_n_423, mul_109_11_n_424, mul_109_11_n_425,
     mul_109_11_n_426, mul_109_11_n_427, mul_109_11_n_428, mul_109_11_n_429,
     mul_109_11_n_430, mul_109_11_n_431, mul_109_11_n_432, mul_109_11_n_433,
     mul_109_11_n_434, mul_109_11_n_435, mul_109_11_n_436, mul_109_11_n_437,
     mul_109_11_n_438, mul_109_11_n_439, mul_109_11_n_440, mul_109_11_n_441,
     mul_109_11_n_442, mul_109_11_n_443, mul_109_11_n_444, mul_109_11_n_445,
     mul_109_11_n_446, mul_109_11_n_447, mul_109_11_n_448, mul_109_11_n_449,
     mul_109_11_n_450, mul_109_11_n_451, mul_109_11_n_452, mul_109_11_n_453,
     mul_109_11_n_454, mul_109_11_n_455, mul_109_11_n_456, mul_109_11_n_457,
     mul_109_11_n_458, mul_109_11_n_459, mul_109_11_n_460, mul_109_11_n_461,
     mul_109_11_n_462, mul_109_11_n_463, mul_109_11_n_464, mul_109_11_n_465,
     mul_109_11_n_466, mul_109_11_n_467, mul_109_11_n_468, mul_109_11_n_469,
     mul_109_11_n_470, mul_109_11_n_471, mul_109_11_n_472, mul_109_11_n_473,
     mul_109_11_n_474, mul_109_11_n_475, mul_109_11_n_476, mul_109_11_n_477,
     mul_109_11_n_478, mul_109_11_n_479, mul_109_11_n_480, mul_109_11_n_481,
     mul_109_11_n_482, mul_109_11_n_483, mul_109_11_n_484, mul_109_11_n_485,
     mul_109_11_n_486, mul_109_11_n_487, mul_109_11_n_488, mul_109_11_n_489,
     mul_109_11_n_490, mul_109_11_n_491, mul_109_11_n_492, mul_109_11_n_493,
     mul_109_11_n_494, mul_109_11_n_495, mul_109_11_n_496, mul_109_11_n_497,
     mul_109_11_n_498, mul_109_11_n_499, mul_109_11_n_500, mul_109_11_n_501,
     mul_109_11_n_502, mul_109_11_n_503, mul_109_11_n_504, mul_109_11_n_505,
     mul_109_11_n_506, mul_109_11_n_507, mul_109_11_n_508, mul_109_11_n_509,
     mul_109_11_n_510, mul_109_11_n_511, mul_109_11_n_512, mul_109_11_n_513,
     mul_109_11_n_514, mul_109_11_n_515, mul_109_11_n_516, mul_109_11_n_517,
     mul_109_11_n_518, mul_109_11_n_519, mul_109_11_n_520, mul_109_11_n_521,
     mul_109_11_n_522, mul_109_11_n_523, mul_109_11_n_524, mul_109_11_n_525,
     mul_109_11_n_526, mul_109_11_n_527, mul_109_11_n_528, mul_109_11_n_529,
     mul_109_11_n_530, mul_109_11_n_531, mul_109_11_n_532, mul_109_11_n_533,
     mul_109_11_n_534, mul_109_11_n_535, mul_109_11_n_536, mul_109_11_n_537,
     mul_109_11_n_538, mul_109_11_n_539, mul_109_11_n_540, mul_109_11_n_541,
     mul_109_11_n_542, mul_109_11_n_543, mul_109_11_n_544, mul_109_11_n_545,
     mul_109_11_n_546, mul_109_11_n_547, mul_109_11_n_548, mul_109_11_n_549,
     mul_109_11_n_550, mul_109_11_n_551, mul_109_11_n_552, mul_109_11_n_553,
     mul_109_11_n_554, mul_109_11_n_555, mul_109_11_n_556, mul_109_11_n_557,
     mul_109_11_n_558, mul_109_11_n_559, mul_109_11_n_560, mul_109_11_n_561,
     mul_109_11_n_562, mul_109_11_n_563, mul_109_11_n_564, mul_109_11_n_565,
     mul_109_11_n_566, mul_109_11_n_567, mul_109_11_n_568, mul_109_11_n_569,
     mul_109_11_n_570, mul_109_11_n_571, mul_109_11_n_572, mul_109_11_n_573,
     mul_109_11_n_574, mul_109_11_n_575, mul_109_11_n_576, mul_109_11_n_577,
     mul_109_11_n_578, mul_109_11_n_579, mul_109_11_n_580, mul_109_11_n_581,
     mul_109_11_n_582, mul_109_11_n_583, mul_109_11_n_584, mul_109_11_n_585,
     mul_109_11_n_586, mul_109_11_n_587, mul_109_11_n_588, mul_109_11_n_589,
     mul_109_11_n_590, mul_109_11_n_591, mul_109_11_n_592, mul_109_11_n_593,
     mul_109_11_n_594, mul_109_11_n_595, mul_109_11_n_596, mul_109_11_n_597,
     mul_109_11_n_598, mul_109_11_n_599, mul_109_11_n_600, mul_109_11_n_601,
     mul_109_11_n_602, mul_109_11_n_603, mul_109_11_n_604, mul_109_11_n_605,
     mul_109_11_n_606, mul_109_11_n_607, mul_109_11_n_608, mul_109_11_n_609,
     mul_109_11_n_610, mul_109_11_n_611, mul_109_11_n_612, mul_109_11_n_613,
     mul_109_11_n_614, mul_109_11_n_615, mul_109_11_n_616, mul_109_11_n_617,
     mul_109_11_n_618, mul_109_11_n_619, mul_109_11_n_620, mul_109_11_n_621,
     mul_109_11_n_622, mul_109_11_n_623, mul_109_11_n_624, mul_109_11_n_625,
     mul_109_11_n_626, mul_109_11_n_627, mul_109_11_n_628, mul_109_11_n_629,
     mul_109_11_n_630, mul_109_11_n_631, mul_109_11_n_632, mul_109_11_n_633,
     mul_109_11_n_634, mul_109_11_n_635, mul_109_11_n_636, mul_109_11_n_637,
     mul_109_11_n_638, mul_109_11_n_639, mul_109_11_n_640, mul_109_11_n_641,
     mul_109_11_n_642, mul_109_11_n_643, mul_109_11_n_644, mul_109_11_n_645,
     mul_109_11_n_646, mul_109_11_n_647, mul_109_11_n_648, mul_109_11_n_649,
     mul_109_11_n_650, mul_109_11_n_651, mul_109_11_n_652, mul_109_11_n_653,
     mul_109_11_n_654, mul_109_11_n_655, mul_109_11_n_656, mul_109_11_n_657,
     mul_109_11_n_658, mul_109_11_n_659, mul_109_11_n_660, mul_109_11_n_661,
     mul_109_11_n_662, mul_109_11_n_663, mul_109_11_n_664, mul_109_11_n_665,
     mul_109_11_n_666, mul_109_11_n_667, mul_109_11_n_668, mul_109_11_n_669,
     mul_109_11_n_670, mul_109_11_n_671, mul_109_11_n_672, mul_109_11_n_673,
     mul_109_11_n_674, mul_109_11_n_675, mul_109_11_n_676, mul_109_11_n_677,
     mul_109_11_n_678, mul_109_11_n_679, mul_109_11_n_680, mul_109_11_n_682,
     mul_109_11_n_683, mul_109_11_n_684, mul_109_11_n_685, mul_109_11_n_686,
     mul_109_11_n_687, mul_109_11_n_688, mul_109_11_n_689, mul_109_11_n_690,
     mul_109_11_n_691, mul_109_11_n_692, mul_109_11_n_693, mul_109_11_n_694,
     mul_109_11_n_695, mul_109_11_n_696, mul_109_11_n_697, mul_109_11_n_698,
     mul_109_11_n_699, mul_109_11_n_700, mul_109_11_n_701, mul_109_11_n_702,
     mul_109_11_n_703, mul_109_11_n_704, mul_109_11_n_705, mul_109_11_n_706,
     mul_109_11_n_707, mul_109_11_n_708, mul_109_11_n_709, mul_109_11_n_710,
     mul_109_11_n_711, mul_109_11_n_712, mul_109_11_n_713, mul_109_11_n_714,
     mul_109_11_n_715, mul_109_11_n_716, mul_109_11_n_717, mul_109_11_n_718,
     mul_109_11_n_719, mul_109_11_n_720, mul_109_11_n_721, mul_109_11_n_722,
     mul_109_11_n_723, mul_109_11_n_724, mul_109_11_n_725, mul_109_11_n_726,
     mul_109_11_n_727, mul_109_11_n_728, mul_109_11_n_729, mul_109_11_n_730,
     mul_109_11_n_731, mul_109_11_n_732, mul_109_11_n_734, mul_109_11_n_735,
     mul_109_11_n_736, mul_109_11_n_737, mul_109_11_n_738, mul_109_11_n_739,
     mul_109_11_n_740, mul_109_11_n_741, mul_109_11_n_742, mul_109_11_n_743,
     mul_109_11_n_744, mul_109_11_n_745, mul_109_11_n_746, mul_109_11_n_747,
     mul_109_11_n_748, mul_109_11_n_749, mul_109_11_n_750, mul_109_11_n_751,
     mul_109_11_n_752, mul_109_11_n_753, mul_109_11_n_754, mul_109_11_n_755,
     mul_109_11_n_756, mul_109_11_n_757, mul_109_11_n_758, mul_109_11_n_759,
     mul_109_11_n_760, mul_109_11_n_761, mul_109_11_n_762, mul_109_11_n_763,
     mul_109_11_n_764, mul_109_11_n_765, mul_109_11_n_766, mul_109_11_n_767,
     mul_109_11_n_768, mul_109_11_n_769, mul_109_11_n_770, mul_109_11_n_771,
     mul_109_11_n_772, mul_109_11_n_773, mul_109_11_n_774, mul_109_11_n_775,
     mul_109_11_n_776, mul_109_11_n_777, mul_109_11_n_778, mul_109_11_n_779,
     mul_109_11_n_780, mul_109_11_n_781, mul_109_11_n_782, mul_109_11_n_783,
     mul_109_11_n_784, mul_109_11_n_785, mul_109_11_n_786, mul_109_11_n_787,
     mul_109_11_n_788, mul_109_11_n_789, mul_109_11_n_790, mul_109_11_n_791,
     mul_109_11_n_792, mul_109_11_n_793, mul_109_11_n_794, mul_109_11_n_795,
     mul_109_11_n_796, mul_109_11_n_797, mul_109_11_n_798, mul_109_11_n_799,
     mul_109_11_n_800, mul_109_11_n_801, mul_109_11_n_802, mul_109_11_n_803,
     mul_109_11_n_805, mul_109_11_n_806, mul_109_11_n_807, mul_109_11_n_808,
     mul_109_11_n_809, mul_109_11_n_810, mul_109_11_n_811, mul_109_11_n_812,
     mul_109_11_n_813, mul_109_11_n_814, mul_109_11_n_815, mul_109_11_n_816,
     mul_109_11_n_817, mul_109_11_n_818, mul_109_11_n_819, mul_109_11_n_820,
     mul_109_11_n_821, mul_109_11_n_822, mul_109_11_n_823, mul_109_11_n_824,
     mul_109_11_n_825, mul_109_11_n_826, mul_109_11_n_827, mul_109_11_n_828,
     mul_109_11_n_829, mul_109_11_n_830, mul_109_11_n_831, mul_109_11_n_832,
     mul_109_11_n_833, mul_109_11_n_834, mul_109_11_n_835, mul_109_11_n_836,
     mul_109_11_n_837, mul_109_11_n_838, mul_109_11_n_839, mul_109_11_n_840,
     mul_109_11_n_841, mul_109_11_n_842, mul_109_11_n_843, mul_109_11_n_844,
     mul_109_11_n_845, mul_109_11_n_846, mul_109_11_n_847, mul_109_11_n_848,
     mul_109_11_n_849, mul_109_11_n_850, mul_109_11_n_851, mul_109_11_n_852,
     mul_109_11_n_853, mul_109_11_n_854, mul_109_11_n_855, mul_109_11_n_856,
     mul_109_11_n_857, mul_109_11_n_858, mul_109_11_n_859, mul_109_11_n_860,
     mul_109_11_n_861, mul_109_11_n_862, mul_109_11_n_863, mul_109_11_n_864,
     mul_109_11_n_865, mul_109_11_n_866, mul_109_11_n_867, mul_109_11_n_868,
     mul_109_11_n_869, mul_109_11_n_870, mul_109_11_n_871, mul_109_11_n_872,
     mul_109_11_n_873, mul_109_11_n_874, mul_109_11_n_875, mul_109_11_n_876,
     mul_109_11_n_877, mul_109_11_n_878, mul_109_11_n_879, mul_109_11_n_880,
     mul_109_11_n_881, mul_109_11_n_882, mul_109_11_n_883, mul_109_11_n_885,
     mul_109_11_n_886, mul_109_11_n_887, mul_109_11_n_888, mul_109_11_n_889,
     mul_109_11_n_890, mul_109_11_n_891, mul_109_11_n_892, mul_109_11_n_893,
     mul_109_11_n_894, mul_109_11_n_895, mul_109_11_n_896, mul_109_11_n_897,
     mul_109_11_n_898, mul_109_11_n_899, mul_109_11_n_900, mul_109_11_n_901,
     mul_109_11_n_902, mul_109_11_n_903, mul_109_11_n_904, mul_109_11_n_905,
     mul_109_11_n_906, mul_109_11_n_907, mul_109_11_n_908, mul_109_11_n_909,
     mul_109_11_n_910, mul_109_11_n_911, mul_109_11_n_912, mul_109_11_n_913,
     mul_109_11_n_914, mul_109_11_n_915, mul_109_11_n_916, mul_109_11_n_917,
     mul_109_11_n_918, mul_109_11_n_919, mul_109_11_n_920, mul_109_11_n_921,
     mul_109_11_n_922, mul_109_11_n_923, mul_109_11_n_924, mul_109_11_n_925,
     mul_109_11_n_926, mul_109_11_n_927, mul_109_11_n_928, mul_109_11_n_929,
     mul_109_11_n_930, mul_109_11_n_931, mul_109_11_n_932, mul_109_11_n_933,
     mul_109_11_n_934, mul_109_11_n_935, mul_109_11_n_936, mul_109_11_n_938,
     mul_109_11_n_939, mul_109_11_n_940, mul_109_11_n_941, mul_109_11_n_942,
     mul_109_11_n_943, mul_109_11_n_944, mul_109_11_n_945, mul_109_11_n_946,
     mul_109_11_n_947, mul_109_11_n_948, mul_109_11_n_949, mul_109_11_n_950,
     mul_109_11_n_951, mul_109_11_n_952, mul_109_11_n_953, mul_109_11_n_954,
     mul_109_11_n_955, mul_109_11_n_956, mul_109_11_n_957, mul_109_11_n_958,
     mul_109_11_n_959, mul_109_11_n_960, mul_109_11_n_961, mul_109_11_n_962,
     mul_109_11_n_963, mul_109_11_n_964, mul_109_11_n_965, mul_109_11_n_966,
     mul_109_11_n_967, mul_109_11_n_968, mul_109_11_n_969, mul_109_11_n_970,
     mul_109_11_n_971, mul_109_11_n_972, mul_109_11_n_973, mul_109_11_n_975,
     mul_109_11_n_976, mul_109_11_n_977, mul_109_11_n_978, mul_109_11_n_979,
     mul_109_11_n_980, mul_109_11_n_981, mul_109_11_n_982, mul_109_11_n_983,
     mul_109_11_n_984, mul_109_11_n_985, mul_109_11_n_986, mul_109_11_n_987,
     mul_109_11_n_988, mul_109_11_n_989, mul_109_11_n_990, mul_109_11_n_991,
     mul_109_11_n_992, mul_109_11_n_993, mul_109_11_n_994, mul_109_11_n_995,
     mul_109_11_n_996, mul_109_11_n_997, mul_109_11_n_998, mul_109_11_n_999,
     mul_109_11_n_1000, mul_109_11_n_1001, mul_109_11_n_1002, mul_109_11_n_1003,
     mul_109_11_n_1004, mul_109_11_n_1005, mul_109_11_n_1006, mul_109_11_n_1007,
     mul_109_11_n_1008, mul_109_11_n_1009, mul_109_11_n_1010, mul_109_11_n_1011,
     mul_109_11_n_1012, mul_109_11_n_1013, mul_109_11_n_1014, mul_109_11_n_1015,
     mul_109_11_n_1016, mul_109_11_n_1017, mul_109_11_n_1018, mul_109_11_n_1019,
     mul_109_11_n_1020, mul_109_11_n_1021, mul_109_11_n_1022, mul_109_11_n_1023,
     mul_109_11_n_1024, mul_109_11_n_1025, mul_109_11_n_1026, mul_109_11_n_1027,
     mul_109_11_n_1028, mul_109_11_n_1029, mul_109_11_n_1030, mul_109_11_n_1031,
     mul_109_11_n_1032, mul_109_11_n_1034, mul_109_11_n_1035, mul_109_11_n_1036,
     mul_109_11_n_1037, mul_109_11_n_1038, mul_109_11_n_1039, mul_109_11_n_1040,
     mul_109_11_n_1041, mul_109_11_n_1042, mul_109_11_n_1043, mul_109_11_n_1044,
     mul_109_11_n_1045, mul_109_11_n_1046, mul_109_11_n_1047, mul_109_11_n_1048,
     mul_109_11_n_1049, mul_109_11_n_1050, mul_109_11_n_1051, mul_109_11_n_1052,
     mul_109_11_n_1053, mul_109_11_n_1054, mul_109_11_n_1055, mul_109_11_n_1056,
     mul_109_11_n_1057, mul_109_11_n_1058, mul_109_11_n_1059, mul_109_11_n_1060,
     mul_109_11_n_1061, mul_109_11_n_1062, mul_109_11_n_1063, mul_109_11_n_1064,
     mul_109_11_n_1065, mul_109_11_n_1066, mul_109_11_n_1067, mul_109_11_n_1068,
     mul_109_11_n_1069, mul_109_11_n_1070, mul_109_11_n_1071, mul_109_11_n_1072,
     mul_109_11_n_1073, mul_109_11_n_1074, mul_109_11_n_1075, mul_109_11_n_1076,
     mul_109_11_n_1077, mul_109_11_n_1078, mul_109_11_n_1079, mul_109_11_n_1080,
     mul_109_11_n_1081, mul_109_11_n_1082, mul_109_11_n_1083, mul_109_11_n_1084,
     mul_109_11_n_1085, mul_109_11_n_1086, mul_109_11_n_1087, mul_109_11_n_1088,
     mul_109_11_n_1089, mul_109_11_n_1090, mul_109_11_n_1092, mul_109_11_n_1093,
     mul_109_11_n_1094, mul_109_11_n_1095, mul_109_11_n_1096, mul_109_11_n_1097,
     mul_109_11_n_1098, mul_109_11_n_1099, mul_109_11_n_1100, mul_109_11_n_1101,
     mul_109_11_n_1102, mul_109_11_n_1103, mul_109_11_n_1104, mul_109_11_n_1105,
     mul_109_11_n_1106, mul_109_11_n_1107, mul_109_11_n_1108, mul_109_11_n_1109,
     mul_109_11_n_1110, mul_109_11_n_1111, mul_109_11_n_1112, mul_109_11_n_1113,
     mul_109_11_n_1114, mul_109_11_n_1115, mul_109_11_n_1116, mul_109_11_n_1117,
     mul_109_11_n_1118, mul_109_11_n_1119, mul_109_11_n_1120, mul_109_11_n_1123,
     mul_109_11_n_1124, mul_109_11_n_1125, mul_109_11_n_1126, mul_109_11_n_1127,
     mul_109_11_n_1128, mul_109_11_n_1129, mul_109_11_n_1130, mul_109_11_n_1131,
     mul_109_11_n_1132, mul_109_11_n_1133, mul_109_11_n_1134, mul_109_11_n_1135,
     mul_109_11_n_1136, mul_109_11_n_1137, mul_109_11_n_1138, mul_109_11_n_1139,
     mul_109_11_n_1140, mul_109_11_n_1141, mul_109_11_n_1142, mul_109_11_n_1143,
     mul_109_11_n_1144, mul_109_11_n_1145, mul_109_11_n_1146, mul_109_11_n_1147,
     mul_109_11_n_1148, mul_109_11_n_1149, mul_109_11_n_1150, mul_109_11_n_1151,
     mul_109_11_n_1154, mul_109_11_n_1155, mul_109_11_n_1156, mul_109_11_n_1157,
     mul_109_11_n_1158, mul_109_11_n_1159, mul_109_11_n_1160, mul_109_11_n_1161,
     mul_109_11_n_1162, mul_109_11_n_1163, mul_109_11_n_1164, mul_109_11_n_1165,
     mul_109_11_n_1166, mul_109_11_n_1167, mul_109_11_n_1168, mul_109_11_n_1169,
     mul_109_11_n_1170, mul_109_11_n_1171, mul_109_11_n_1172, mul_109_11_n_1173,
     mul_109_11_n_1174, mul_109_11_n_1175, mul_109_11_n_1176, mul_109_11_n_1177,
     mul_109_11_n_1178, mul_109_11_n_1179, mul_109_11_n_1182, mul_109_11_n_1183,
     mul_109_11_n_1184, mul_109_11_n_1185, mul_109_11_n_1186, mul_109_11_n_1187,
     mul_109_11_n_1188, mul_109_11_n_1189, mul_109_11_n_1190, mul_109_11_n_1191,
     mul_109_11_n_1192, mul_109_11_n_1193, mul_109_11_n_1194, mul_109_11_n_1195,
     mul_109_11_n_1196, mul_109_11_n_1197, mul_109_11_n_1198, mul_109_11_n_1199,
     mul_109_11_n_1200, mul_109_11_n_1201, mul_109_11_n_1202, mul_109_11_n_1203,
     mul_109_11_n_1205, mul_109_11_n_1206, mul_109_11_n_1207, mul_109_11_n_1208,
     mul_109_11_n_1209, mul_109_11_n_1210, mul_109_11_n_1211, mul_109_11_n_1212,
     mul_109_11_n_1213, mul_109_11_n_1214, mul_109_11_n_1215, mul_109_11_n_1216,
     mul_109_11_n_1217, mul_109_11_n_1218, mul_109_11_n_1219, mul_109_11_n_1220,
     mul_109_11_n_1221, mul_109_11_n_1222, mul_109_11_n_1223, mul_109_11_n_1224,
     mul_109_11_n_1225, mul_109_11_n_1226, mul_109_11_n_1227, mul_109_11_n_1228,
     mul_109_11_n_1229, mul_109_11_n_1230, mul_109_11_n_1231, mul_109_11_n_1232,
     mul_109_11_n_1233, mul_109_11_n_1234, mul_109_11_n_1235, mul_109_11_n_1236,
     mul_109_11_n_1237, mul_109_11_n_1238, mul_109_11_n_1239, mul_109_11_n_1240,
     mul_109_11_n_1241, mul_109_11_n_1242, mul_109_11_n_1243, mul_109_11_n_1244,
     mul_109_11_n_1245, mul_109_11_n_1246, mul_109_11_n_1247, mul_109_11_n_1248,
     mul_109_11_n_1249, mul_109_11_n_1250, mul_109_11_n_1251, mul_109_11_n_1252,
     mul_109_11_n_1253, mul_109_11_n_1254, mul_109_11_n_1255, mul_109_11_n_1256,
     mul_109_11_n_1257, mul_109_11_n_1258, mul_109_11_n_1259, mul_109_11_n_1260,
     mul_109_11_n_1261, mul_109_11_n_1264, mul_109_11_n_1265, mul_109_11_n_1266,
     mul_109_11_n_1267, mul_109_11_n_1268, mul_109_11_n_1269, mul_109_11_n_1270,
     mul_109_11_n_1271, mul_109_11_n_1273, mul_109_11_n_1274, mul_109_11_n_1275,
     mul_109_11_n_1276, mul_109_11_n_1277, mul_109_11_n_1278, mul_109_11_n_1279,
     mul_109_11_n_1280, mul_109_11_n_1282, mul_109_11_n_1285, mul_109_11_n_1286,
     mul_109_11_n_1287, mul_109_11_n_1290, mul_109_11_n_1291, mul_109_11_n_1292,
     mul_109_11_n_1294, mul_109_11_n_1296, mul_109_11_n_1297, mul_109_11_n_1300,
     mul_109_11_n_1301, mul_109_11_n_1303, mul_109_11_n_1304, n_0, n_1, n_2, n_3,
     n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15, n_16,
     n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26, n_27, n_28,
     n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39, n_40,
     n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50, n_51, n_52,
     n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64,
     n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76,
     n_77, n_78, n_79, n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88,
     n_89, n_90, n_91, n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100,
     n_101, n_102, n_103, n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111,
     n_112, n_113, n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122,
     n_123, n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133,
     n_134, n_135, n_136, n_137, n_138, n_139, n_140, n_141, n_142, n_143, n_144,
     n_145, n_146, n_147, n_148, n_149, n_150, n_151, n_152, n_153, n_154, n_155,
     n_156, n_157, n_158, n_159, n_160, n_161, n_162, n_163, n_164, n_165, n_166,
     n_167, n_168, n_169, n_170, n_171, n_172, n_173, n_174, n_175, n_176, n_177,
     n_178, n_179, n_180, n_181, n_182, n_183, n_184, n_185, n_186, n_187, n_188,
     n_189, n_190, n_191, n_192, n_193, n_194, n_195, n_196, n_197, n_198, n_199,
     n_200, n_201, n_202, n_203, n_204, n_205, n_206, n_207, n_208, n_209, n_210,
     n_211, n_212, n_213, n_214, n_215, n_216, n_217, n_218, n_219, n_220, n_221,
     n_222, n_223, n_224, n_225, n_226, n_227, n_228, n_229, n_230, n_231, n_232,
     n_233, n_234, n_235, n_236, n_237, n_238, n_239, n_240, n_241, n_242, n_243,
     n_244, n_245, n_246, n_247, n_248, n_249, n_250, n_251, n_252, n_253, n_254,
     n_255, n_256, n_257, n_258, n_259, n_260, n_261, n_262, n_263, n_264, n_265,
     n_266, n_267, n_268, n_269, n_270, n_271, n_272, n_273, n_274, n_275, n_276,
     n_277, n_310, n_311, n_312, n_313, n_314, n_315, n_316, n_317, n_318, n_319,
     n_320, n_321, n_322, n_323, n_324, n_325, n_326, n_327, n_328, n_329, n_330,
     n_331, n_332, n_333, n_334, n_335, n_336, n_337, n_338, n_339, n_340, n_341,
     n_342, n_343, n_344, n_345, n_346, n_347, n_348, n_349, n_350, n_351, n_352,
     n_353, n_354, n_355, n_356, n_357, n_358, n_359, n_360, n_361, n_362, n_363,
     n_364, n_365, n_366, n_367, n_368, n_369, n_370, n_371, n_372, n_373, n_374,
     n_375, n_376, n_377, n_378, n_379, n_380, n_381, n_382, n_383, n_384, n_385,
     n_386, n_387, n_388, n_389, n_390, n_391, n_392, n_393, n_394, n_395, n_396,
     n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404, n_405, n_406, n_407,
     n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415, n_416, n_417, n_418,
     n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426, n_427, n_428, n_429,
     n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437, n_438, n_439, n_440,
     n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448, n_449, n_450, n_451,
     n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459, n_460, n_461, n_462,
     n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470, n_471, n_472, n_473,
     n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481, n_482, n_483, n_484,
     n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492, n_493, n_494, n_495,
     n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503, n_504, n_505, n_506,
     n_507, n_508, n_509, n_510, n_511, n_512, n_513, n_514, n_515, n_516, n_517,
     n_518, n_519, n_520, n_521, n_522, n_523, n_524, n_525, n_526, n_527, n_528,
     n_529, n_530, n_531, n_532, n_533, n_534, n_535, n_536, n_537, n_538, n_539,
     n_540, n_541, n_542, n_543, n_544, n_545, n_546, n_547, n_548, n_549, n_550,
     n_551, n_552, n_553, n_554, n_555, n_556, n_557, n_558, n_559, n_560, n_561,
     n_562, n_563, n_564, n_565, n_566, n_567, n_568, n_569, n_570, n_571, n_572,
     n_573, n_574, n_575, n_576, n_577, n_578, n_579, n_580, n_581, n_582, n_583,
     n_584, n_585, n_586, n_587, n_588, n_589, n_590, n_591, n_592, n_593, n_594,
     n_595, n_596, n_597, n_598, n_599, n_600, n_601, n_602, n_603, n_604, n_605,
     n_606, n_607, n_608, n_609, n_610, n_611, n_612, n_613, n_614, n_615, n_616,
     n_617, n_618, n_619, clk, stall, n_654, n_655, n_656, n_657, n_658, n_659,
     n_660, n_661, n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_669, n_670,
     n_671, n_672, n_673, n_674, n_675, n_676, n_677, n_678, n_679, n_680, n_681,
     n_682, n_683, n_684, n_685, n_686, n_687, n_688, n_689, n_690, n_691, n_692,
     n_693, n_694, n_695, n_696, n_697, n_698, n_699, n_700, n_701, n_702, n_703,
     n_704, n_705, n_706, n_707, n_708, n_709, n_710, n_711, n_712, n_713, n_714,
     n_715, n_716, n_717, n_718, n_719, n_720, n_721, n_722, n_723, n_724, n_725,
     n_726, n_727, n_728, n_729, n_730, n_731, n_732, n_733, n_734, n_735, n_736,
     n_737, n_738, n_739, n_740, n_741, n_742, n_743, n_744, n_745, n_746, n_747,
     n_748, n_749, n_750, n_751, n_752, n_753, n_754, n_755, n_756, n_757, n_758,
     n_759, n_760, n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768, n_769,
     n_770, n_771, n_772, n_773, n_774, n_775, n_776, n_777, n_778, n_779, n_780,
     n_781, n_782, n_783, n_784, n_785, n_786, n_787, n_788, n_789, n_790, n_791,
     n_792, n_793, n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801, n_802,
     n_803, n_804, n_805, n_806, n_807, n_808, n_809, n_810, n_811, n_812, n_813,
     n_814, n_815, n_816, n_817, n_818, n_819, n_820, n_821, n_822, n_823, n_824,
     n_825, n_826, n_827, n_828, n_829, n_830, n_831, n_832, n_833, n_834, n_835,
     n_836, n_837, n_838, n_839, n_840, n_841, n_842, n_843, n_844, n_845, n_846,
     n_847, n_848, n_849, n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857,
     n_858, n_859, n_860, n_861, n_862, n_863, n_864, n_865, n_866, n_867, n_868,
     n_869, n_870, n_871, n_872, n_873, n_874, n_875, n_876, n_877, n_878, n_879,
     n_880, n_881, n_882, n_883, n_884, n_885, n_886, n_887, n_888, n_889, n_890,
     n_891, n_892, n_893, n_894, n_895, n_896, n_897, n_898, n_899, n_900, n_901,
     n_902, n_903, n_904, n_905, n_906, n_907, n_908, n_909, n_910, n_911, n_913,
     n_914, n_915, n_916, n_917, n_918, n_919, n_920, n_921, n_922, n_923, n_924,
     n_925, n_926, n_927, n_928, n_929, n_930, n_931, n_932, n_933, n_934, n_935,
     n_936, n_937, n_938, n_939, n_940, n_941, n_942, n_943, n_944, n_945, n_946,
     n_947, n_948, n_949, n_950, n_951, n_952, n_953, n_954, n_955, n_956, n_957,
     n_958, n_959, n_960, n_961, n_962, n_963, n_964, n_965, n_966, n_967, n_968,
     n_969, n_970, n_971, n_972, n_973, n_974, n_975, n_976, n_977, n_978, n_979,
     n_980, n_981, n_982, n_983, n_984, n_985, n_986, n_987, n_988, n_989, n_990,
     n_991, n_992, n_993, n_994, n_995, n_996, n_997, n_998, n_999, n_1000,
     n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007, n_1008, n_1009,
     n_1010, n_1011, n_1012, n_1013, n_1014, n_1015, n_1016, n_1017, n_1018,
     n_1019, n_1020, n_1021, n_1022, n_1023, n_1024, n_1025, n_1026, n_1027,
     n_1028, n_1029, n_1030, n_1031, n_1032, n_1033, n_1034, n_1035, n_1036,
     n_1037, n_1038, n_1039, n_1040, n_1041, n_1042, n_1043, n_1044, n_1045,
     n_1046, n_1047, n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054,
     n_1055, n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063,
     n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071, n_1072,
     n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079, n_1080, n_1081,
     n_1082, n_1083, n_1084, n_1085, n_1086, n_1087, n_1088, n_1089, n_1090,
     n_1091, n_1092, n_1093, n_1094, n_1095, n_1096, n_1097, n_1098, n_1099,
     n_1100, n_1101, n_1102, n_1103, n_1104, n_1105, n_1106, n_1107, n_1108,
     n_1109, n_1110, n_1111, n_1112, n_1113, n_1114, n_1115, n_1116, n_1117,
     n_1118, n_1119, n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126,
     n_1127, n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135,
     n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143, n_1144,
     n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151, n_1152, n_1153,
     n_1154, n_1155, n_1156, n_1157, n_1158, n_1159, n_1160, n_1161, n_1162,
     n_1163, n_1164, n_1165, n_1166, n_1167, n_1168, n_1169, n_1170, n_1171,
     n_1172, n_1173, n_1174, n_1175, n_1176, n_1177, n_1178, n_1179, n_1180,
     n_1181, n_1182, n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1189,
     n_1190, n_1191, n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198,
     n_1199, n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207,
     n_1208, n_1209, n_1274, n_1275, n_1276, n_1277, n_1278, n_1279, n_1280,
     n_1282, n_1283, n_1284, n_1285, n_1286, n_1287, n_1292, n_1294, n_1295,
     n_1296, n_1297, n_1298, n_1299, n_1300, n_1301, n_1302, n_1303, n_1304,
     n_1306, n_1309, n_1310, n_1311, n_1312, n_1313, n_1314, n_1315, n_1316,
     n_1317, n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325,
     n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333, n_1334,
     n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341, n_1344, n_1346,
     n_1347, n_1348, n_1349, n_1350, n_1351, n_1352, n_1353, n_1354, n_1355,
     n_1356, n_1357, n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364,
     n_1365, n_1366, n_1367, n_1368, n_1369, n_1370, n_1371, n_1372, n_1373,
     n_1374, n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382,
     n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390, n_1391,
     n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398, n_1399, n_1400,
     n_1401, n_1402, n_1403, n_1404, n_1405, n_1406, n_1407, n_1408, n_1409,
     n_1410, n_1411, n_1412, n_1413, n_1414, n_1415, n_1416, n_1417, n_1418,
     n_1419, n_1420, n_1421, n_1422, n_1423, n_1424, n_1425, n_1426, n_1427,
     n_1428, n_1429, n_1430, n_1431, n_1432, n_1433, n_1434, n_1435, n_1436,
     n_1437, n_1438, n_1439, n_1440, n_1441, n_1442, n_1443, n_1444, n_1445,
     n_1446, n_1447, n_1448, n_1449, n_1450, n_1451, n_1452, n_1453, n_1454,
     n_1455, n_1456, n_1457, n_1458, n_1459, n_1460, n_1461, n_1462, n_1463,
     n_1464, n_1465, n_1466, n_1467, n_1468, n_1470, n_1471, n_1472, n_1473,
     n_1474, n_1476, n_1477, n_1478, n_1479, n_1480, n_1481, n_1482, n_1483,
     n_1484, n_1485, n_1486, n_1487, n_1488, n_1489, n_1490, n_1491, n_1492,
     n_1493, n_1494, n_1495, n_1496, n_1497, n_1498, n_1499, n_1500, n_1501,
     n_1502, n_1503, n_1504, n_1505, n_1506, n_1507, n_1508, n_1509, n_1510,
     n_1511, n_1512, n_1513, n_1514, n_1515, n_1516, n_1517, n_1518, n_1519,
     n_1520, n_1521, n_1522, n_1523, n_1524, n_1525, n_1526, n_1527, n_1528,
     n_1529, n_1530, n_1531, n_1532, n_1533, n_1534;
 reg retime_s1_1_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s1_1_reg_reg_N30 <= n_567;
 assign n_0 = retime_s1_1_reg_reg_N30;
 reg retime_s1_2_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_2_reg_reg_N30 <= {in5[2]};
 assign n_2 = retime_s1_2_reg_reg_N30;
 reg retime_s1_3_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_3_reg_reg_N30 <= csa_tree_add_86_2_n_25;
 assign n_8 = retime_s1_3_reg_reg_N30;
 reg retime_s1_4_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_4_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_46;
 assign n_78 = retime_s1_4_reg_reg_N30;
 reg retime_s1_5_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s1_5_reg_reg_N30 <= n_524;
 assign n_89 = retime_s1_5_reg_reg_N30;
 reg retime_s1_6_reg_reg_N30;
 always @(posedge clk)
         retime_s1_6_reg_reg_N30 <= n_510;
 assign n_91 = retime_s1_6_reg_reg_N30;
 reg retime_s1_7_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_7_reg_reg_N30 <= n_507;
 assign n_93 = retime_s1_7_reg_reg_N30;
 reg retime_s1_8_reg_reg_N30;
 always @(posedge clk)
         retime_s1_8_reg_reg_N30 <= n_501;
 assign n_94 = retime_s1_8_reg_reg_N30;
 reg retime_s1_9_reg_reg_N30;
 always @(posedge clk)
         retime_s1_9_reg_reg_N30 <= n_713;
 assign csa_tree_add_106_2_groupi_n_227 = retime_s1_9_reg_reg_N30;
 reg retime_s1_10_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_10_reg_reg_N30 <= n_980;
 assign n_103 = retime_s1_10_reg_reg_N30;
 reg retime_s1_11_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_11_reg_reg_N30 <= n_1444;
 assign n_104 = retime_s1_11_reg_reg_N30;
 reg retime_s1_12_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s1_12_reg_reg_N30 <= n_195;
 assign n_105 = retime_s1_12_reg_reg_N30;
 reg retime_s1_13_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_13_reg_reg_N30 <= n_1154;
 assign n_107 = retime_s1_13_reg_reg_N30;
 reg retime_s1_14_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_14_reg_reg_N30 <= n_688;
 assign n_108 = retime_s1_14_reg_reg_N30;
 reg retime_s1_15_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_15_reg_reg_N30 <= n_779;
 assign n_109 = retime_s1_15_reg_reg_N30;
 reg retime_s1_16_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_16_reg_reg_N30 <= n_970;
 assign n_110 = retime_s1_16_reg_reg_N30;
 reg retime_s1_17_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_17_reg_reg_N30 <= n_969;
 assign n_111 = retime_s1_17_reg_reg_N30;
 reg retime_s1_18_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_18_reg_reg_N30 <= n_927;
 assign n_112 = retime_s1_18_reg_reg_N30;
 reg retime_s1_19_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_19_reg_reg_N30 <= {in5[4]};
 assign n_113 = retime_s1_19_reg_reg_N30;
 reg retime_s1_20_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_20_reg_reg_N30 <= csa_tree_add_86_2_n_3;
 assign n_114 = retime_s1_20_reg_reg_N30;
 reg retime_s1_21_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_21_reg_reg_N30 <= n_964;
 assign n_115 = retime_s1_21_reg_reg_N30;
 reg retime_s1_22_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_22_reg_reg_N30 <= n_963;
 assign n_116 = retime_s1_22_reg_reg_N30;
 reg retime_s1_23_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_23_reg_reg_N30 <= n_530;
 assign n_117 = retime_s1_23_reg_reg_N30;
 reg retime_s1_24_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_24_reg_reg_N30 <= n_519;
 assign n_118 = retime_s1_24_reg_reg_N30;
 reg retime_s1_25_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_25_reg_reg_N30 <= n_515;
 assign n_119 = retime_s1_25_reg_reg_N30;
 reg retime_s1_26_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_26_reg_reg_N30 <= n_939;
 assign n_120 = retime_s1_26_reg_reg_N30;
 reg retime_s1_27_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_27_reg_reg_N30 <= n_1002;
 assign n_121 = retime_s1_27_reg_reg_N30;
 reg retime_s1_28_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_28_reg_reg_N30 <= n_1001;
 assign n_122 = retime_s1_28_reg_reg_N30;
 reg retime_s1_29_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_29_reg_reg_N30 <= n_707;
 assign n_123 = retime_s1_29_reg_reg_N30;
 reg retime_s1_30_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_30_reg_reg_N30 <= n_706;
 assign n_124 = retime_s1_30_reg_reg_N30;
 reg retime_s1_31_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_31_reg_reg_N30 <= n_583;
 assign n_125 = retime_s1_31_reg_reg_N30;
 reg retime_s1_32_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_32_reg_reg_N30 <= n_582;
 assign n_126 = retime_s1_32_reg_reg_N30;
 reg retime_s1_33_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_33_reg_reg_N30 <= n_1000;
 assign n_127 = retime_s1_33_reg_reg_N30;
 reg retime_s1_34_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_34_reg_reg_N30 <= n_999;
 assign n_128 = retime_s1_34_reg_reg_N30;
 reg retime_s1_35_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_35_reg_reg_N30 <= n_1464;
 assign n_129 = retime_s1_35_reg_reg_N30;
 reg retime_s1_36_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_36_reg_reg_N30 <= n_277;
 assign n_130 = retime_s1_36_reg_reg_N30;
 reg retime_s1_37_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s1_37_reg_reg_N30 <= n_1459;
 assign n_131 = retime_s1_37_reg_reg_N30;
 reg retime_s1_38_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_38_reg_reg_N30 <= n_613;
 assign n_132 = retime_s1_38_reg_reg_N30;
 reg retime_s1_39_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_39_reg_reg_N30 <= n_998;
 assign n_133 = retime_s1_39_reg_reg_N30;
 reg retime_s1_40_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_40_reg_reg_N30 <= n_997;
 assign n_134 = retime_s1_40_reg_reg_N30;
 reg retime_s1_41_reg_reg_N30;
 always @(posedge clk)
         retime_s1_41_reg_reg_N30 <= n_1054;
 assign csa_tree_mul_77_11_groupi_n_594 = retime_s1_41_reg_reg_N30;
 reg retime_s1_42_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_42_reg_reg_N30 <= n_1465;
 assign n_137 = retime_s1_42_reg_reg_N30;
 reg retime_s1_43_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_43_reg_reg_N30 <= n_928;
 assign n_138 = retime_s1_43_reg_reg_N30;
 reg retime_s1_44_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_44_reg_reg_N30 <= n_198;
 assign n_139 = retime_s1_44_reg_reg_N30;
 reg retime_s1_45_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_45_reg_reg_N30 <= n_197;
 assign n_140 = retime_s1_45_reg_reg_N30;
 reg retime_s1_46_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_46_reg_reg_N30 <= n_968;
 assign n_141 = retime_s1_46_reg_reg_N30;
 reg retime_s1_47_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_47_reg_reg_N30 <= n_984;
 assign n_142 = retime_s1_47_reg_reg_N30;
 reg retime_s1_48_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_48_reg_reg_N30 <= n_983;
 assign n_143 = retime_s1_48_reg_reg_N30;
 reg retime_s1_49_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_49_reg_reg_N30 <= n_670;
 assign n_144 = retime_s1_49_reg_reg_N30;
 reg retime_s1_50_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_50_reg_reg_N30 <= n_669;
 assign n_145 = retime_s1_50_reg_reg_N30;
 reg retime_s1_51_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_51_reg_reg_N30 <= n_946;
 assign n_146 = retime_s1_51_reg_reg_N30;
 reg retime_s1_52_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_52_reg_reg_N30 <= n_945;
 assign n_147 = retime_s1_52_reg_reg_N30;
 reg retime_s1_53_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_53_reg_reg_N30 <= n_1463;
 assign n_148 = retime_s1_53_reg_reg_N30;
 reg retime_s1_54_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_54_reg_reg_N30 <= n_535;
 assign n_149 = retime_s1_54_reg_reg_N30;
 reg retime_s1_55_reg_reg_N30;
 always @(posedge clk)
         retime_s1_55_reg_reg_N30 <= n_685;
 assign n_150 = retime_s1_55_reg_reg_N30;
 reg retime_s1_56_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s1_56_reg_reg_N30 <= n_793;
 assign n_151 = retime_s1_56_reg_reg_N30;
 reg retime_s1_57_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_57_reg_reg_N30 <= n_1384;
 assign n_152 = retime_s1_57_reg_reg_N30;
 reg retime_s1_58_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_58_reg_reg_N30 <= n_256;
 assign n_153 = retime_s1_58_reg_reg_N30;
 reg retime_s1_59_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_59_reg_reg_N30 <= n_249;
 assign n_154 = retime_s1_59_reg_reg_N30;
 reg retime_s1_60_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_60_reg_reg_N30 <= n_994;
 assign n_155 = retime_s1_60_reg_reg_N30;
 reg retime_s1_61_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_61_reg_reg_N30 <= n_697;
 assign n_156 = retime_s1_61_reg_reg_N30;
 reg retime_s1_62_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_62_reg_reg_N30 <= n_696;
 assign n_157 = retime_s1_62_reg_reg_N30;
 reg retime_s1_63_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_63_reg_reg_N30 <= n_982;
 assign n_158 = retime_s1_63_reg_reg_N30;
 reg retime_s1_64_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_64_reg_reg_N30 <= n_981;
 assign n_159 = retime_s1_64_reg_reg_N30;
 reg retime_s1_65_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_65_reg_reg_N30 <= n_1431;
 assign n_160 = retime_s1_65_reg_reg_N30;
 reg retime_s1_66_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_66_reg_reg_N30 <= n_938;
 assign n_161 = retime_s1_66_reg_reg_N30;
 reg retime_s1_67_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_67_reg_reg_N30 <= n_200;
 assign n_162 = retime_s1_67_reg_reg_N30;
 reg retime_s1_68_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_68_reg_reg_N30 <= n_199;
 assign n_163 = retime_s1_68_reg_reg_N30;
 reg retime_s1_69_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_69_reg_reg_N30 <= n_931;
 assign n_164 = retime_s1_69_reg_reg_N30;
 reg retime_s1_70_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_70_reg_reg_N30 <= n_930;
 assign n_165 = retime_s1_70_reg_reg_N30;
 reg retime_s1_71_reg_reg_N30;
 always @(posedge clk)
         retime_s1_71_reg_reg_N30 <= n_785;
 assign n_166 = retime_s1_71_reg_reg_N30;
 reg retime_s1_72_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_72_reg_reg_N30 <= n_935;
 assign n_167 = retime_s1_72_reg_reg_N30;
 reg retime_s1_73_reg_reg_N30;
 always @(posedge clk)
         retime_s1_73_reg_reg_N30 <= n_614;
 assign csa_tree_add_106_2_groupi_n_229 = retime_s1_73_reg_reg_N30;
 reg retime_s1_74_reg_reg_N30;
 always @(posedge clk)
         retime_s1_74_reg_reg_N30 <= n_682;
 assign csa_tree_add_106_2_groupi_n_335 = retime_s1_74_reg_reg_N30;
 reg retime_s1_75_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_75_reg_reg_N30 <= n_966;
 assign n_168 = retime_s1_75_reg_reg_N30;
 reg retime_s1_76_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_76_reg_reg_N30 <= n_965;
 assign n_169 = retime_s1_76_reg_reg_N30;
 reg retime_s1_77_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_77_reg_reg_N30 <= n_1339;
 assign n_170 = retime_s1_77_reg_reg_N30;
 reg retime_s1_78_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s1_78_reg_reg_N30 <= n_702;
 assign n_171 = retime_s1_78_reg_reg_N30;
 reg retime_s1_79_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_79_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_113;
 assign n_312 = retime_s1_79_reg_reg_N30;
 reg retime_s1_80_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_80_reg_reg_N30 <= n_972;
 assign n_313 = retime_s1_80_reg_reg_N30;
 reg retime_s1_81_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_81_reg_reg_N30 <= n_971;
 assign n_314 = retime_s1_81_reg_reg_N30;
 reg retime_s1_82_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_82_reg_reg_N30 <= n_666;
 assign n_315 = retime_s1_82_reg_reg_N30;
 reg retime_s1_83_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_83_reg_reg_N30 <= n_665;
 assign n_316 = retime_s1_83_reg_reg_N30;
 reg retime_s1_84_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_84_reg_reg_N30 <= n_710;
 assign n_317 = retime_s1_84_reg_reg_N30;
 reg retime_s1_85_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_85_reg_reg_N30 <= n_675;
 assign n_318 = retime_s1_85_reg_reg_N30;
 reg retime_s1_86_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_86_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_233;
 assign n_319 = retime_s1_86_reg_reg_N30;
 reg retime_s1_87_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_87_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_177;
 assign n_320 = retime_s1_87_reg_reg_N30;
 reg retime_s1_88_reg_reg_N30;
 always @(posedge clk)
         retime_s1_88_reg_reg_N30 <= n_784;
 assign n_321 = retime_s1_88_reg_reg_N30;
 reg retime_s1_89_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_89_reg_reg_N30 <= n_1440;
 assign n_322 = retime_s1_89_reg_reg_N30;
 reg retime_s1_90_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_90_reg_reg_N30 <= n_950;
 assign n_323 = retime_s1_90_reg_reg_N30;
 reg retime_s1_91_reg_reg_N30;
 always @(posedge clk)
         retime_s1_91_reg_reg_N30 <= n_615;
 assign n_324 = retime_s1_91_reg_reg_N30;
 reg retime_s1_92_reg_reg_N30;
 always @(posedge clk)
         retime_s1_92_reg_reg_N30 <= n_616;
 assign n_325 = retime_s1_92_reg_reg_N30;
 reg retime_s1_93_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_93_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_119;
 assign n_326 = retime_s1_93_reg_reg_N30;
 reg retime_s1_94_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_94_reg_reg_N30 <= n_1498;
 assign n_327 = retime_s1_94_reg_reg_N30;
 reg retime_s1_95_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_95_reg_reg_N30 <= n_564;
 assign n_328 = retime_s1_95_reg_reg_N30;
 reg retime_s1_96_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_96_reg_reg_N30 <= n_563;
 assign n_329 = retime_s1_96_reg_reg_N30;
 reg retime_s1_97_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_97_reg_reg_N30 <= n_990;
 assign n_330 = retime_s1_97_reg_reg_N30;
 reg retime_s1_98_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_98_reg_reg_N30 <= n_961;
 assign n_331 = retime_s1_98_reg_reg_N30;
 reg retime_s1_99_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_99_reg_reg_N30 <= n_960;
 assign n_332 = retime_s1_99_reg_reg_N30;
 reg retime_s1_100_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_100_reg_reg_N30 <= n_953;
 assign n_333 = retime_s1_100_reg_reg_N30;
 reg retime_s1_101_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_101_reg_reg_N30 <= n_952;
 assign n_334 = retime_s1_101_reg_reg_N30;
 reg retime_s1_102_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_102_reg_reg_N30 <= n_992;
 assign n_335 = retime_s1_102_reg_reg_N30;
 reg retime_s1_103_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_103_reg_reg_N30 <= n_991;
 assign n_336 = retime_s1_103_reg_reg_N30;
 reg retime_s1_104_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_104_reg_reg_N30 <= n_948;
 assign n_337 = retime_s1_104_reg_reg_N30;
 reg retime_s1_105_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_105_reg_reg_N30 <= n_947;
 assign n_338 = retime_s1_105_reg_reg_N30;
 reg retime_s1_106_reg_reg_N30;
 always @(posedge clk)
         retime_s1_106_reg_reg_N30 <= n_1159;
 assign n_339 = retime_s1_106_reg_reg_N30;
 reg retime_s1_107_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_107_reg_reg_N30 <= n_1466;
 assign n_340 = retime_s1_107_reg_reg_N30;
 reg retime_s1_108_reg_reg_N30;
 always @(posedge clk)
         retime_s1_108_reg_reg_N30 <= n_226;
 assign n_341 = retime_s1_108_reg_reg_N30;
 reg retime_s1_109_reg_reg_N30;
 always @(posedge clk)
         retime_s1_109_reg_reg_N30 <= n_1055;
 assign n_342 = retime_s1_109_reg_reg_N30;
 reg retime_s1_110_reg_reg_N30;
 always @(posedge clk)
         retime_s1_110_reg_reg_N30 <= n_591;
 assign n_343 = retime_s1_110_reg_reg_N30;
 reg retime_s1_111_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_111_reg_reg_N30 <= n_1005;
 assign n_344 = retime_s1_111_reg_reg_N30;
 reg retime_s1_112_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_112_reg_reg_N30 <= n_1004;
 assign n_345 = retime_s1_112_reg_reg_N30;
 reg retime_s1_113_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_113_reg_reg_N30 <= n_956;
 assign n_346 = retime_s1_113_reg_reg_N30;
 reg retime_s1_114_reg_reg_N30;
 always @(posedge clk)
         retime_s1_114_reg_reg_N30 <= n_593;
 assign n_347 = retime_s1_114_reg_reg_N30;
 reg retime_s1_115_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_115_reg_reg_N30 <= n_179;
 assign n_348 = retime_s1_115_reg_reg_N30;
 reg retime_s1_116_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_116_reg_reg_N30 <= n_1344;
 assign n_349 = retime_s1_116_reg_reg_N30;
 reg retime_s1_117_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_117_reg_reg_N30 <= n_1496;
 assign n_350 = retime_s1_117_reg_reg_N30;
 reg retime_s1_118_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_118_reg_reg_N30 <= n_1498;
 assign n_351 = retime_s1_118_reg_reg_N30;
 reg retime_s1_119_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_119_reg_reg_N30 <= n_663;
 assign n_352 = retime_s1_119_reg_reg_N30;
 reg retime_s1_120_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_120_reg_reg_N30 <= n_662;
 assign n_353 = retime_s1_120_reg_reg_N30;
 reg retime_s1_121_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_121_reg_reg_N30 <= n_701;
 assign n_354 = retime_s1_121_reg_reg_N30;
 reg retime_s1_122_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_122_reg_reg_N30 <= n_1495;
 assign n_355 = retime_s1_122_reg_reg_N30;
 reg retime_s1_123_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_123_reg_reg_N30 <= n_955;
 assign n_356 = retime_s1_123_reg_reg_N30;
 reg retime_s1_124_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_124_reg_reg_N30 <= n_1497;
 assign n_357 = retime_s1_124_reg_reg_N30;
 reg retime_s1_125_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_125_reg_reg_N30 <= n_1346;
 assign n_358 = retime_s1_125_reg_reg_N30;
 reg retime_s1_126_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_126_reg_reg_N30 <= n_1346;
 assign n_359 = retime_s1_126_reg_reg_N30;
 reg retime_s1_127_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_127_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_248;
 assign n_360 = retime_s1_127_reg_reg_N30;
 reg retime_s1_128_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_128_reg_reg_N30 <= n_943;
 assign n_361 = retime_s1_128_reg_reg_N30;
 reg retime_s1_129_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_129_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_21;
 assign n_363 = retime_s1_129_reg_reg_N30;
 reg retime_s1_130_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_130_reg_reg_N30 <= n_560;
 assign n_364 = retime_s1_130_reg_reg_N30;
 reg retime_s1_131_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_131_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_48;
 assign n_365 = retime_s1_131_reg_reg_N30;
 reg retime_s1_132_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_132_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_170;
 assign n_366 = retime_s1_132_reg_reg_N30;
 reg retime_s1_133_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_133_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_15;
 assign n_367 = retime_s1_133_reg_reg_N30;
 reg retime_s1_134_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_134_reg_reg_N30 <= n_932;
 assign n_368 = retime_s1_134_reg_reg_N30;
 reg retime_s1_135_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_135_reg_reg_N30 <= n_1171;
 assign n_369 = retime_s1_135_reg_reg_N30;
 reg retime_s1_136_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_136_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_224;
 assign n_371 = retime_s1_136_reg_reg_N30;
 reg retime_s1_137_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_137_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_262;
 assign n_372 = retime_s1_137_reg_reg_N30;
 reg retime_s1_138_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s1_138_reg_reg_N30 <= n_693;
 assign n_373 = retime_s1_138_reg_reg_N30;
 reg retime_s1_139_reg_reg_N30;
 always @(posedge clk)
         retime_s1_139_reg_reg_N30 <= n_221;
 assign n_374 = retime_s1_139_reg_reg_N30;
 reg retime_s1_140_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_140_reg_reg_N30 <= n_1340;
 assign n_375 = retime_s1_140_reg_reg_N30;
 reg retime_s1_141_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_141_reg_reg_N30 <= csa_tree_add_86_2_n_27;
 assign n_376 = retime_s1_141_reg_reg_N30;
 reg retime_s1_142_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_142_reg_reg_N30 <= n_1341;
 assign n_377 = retime_s1_142_reg_reg_N30;
 reg retime_s1_143_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_143_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_222;
 assign n_378 = retime_s1_143_reg_reg_N30;
 reg retime_s1_144_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_144_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_3;
 assign n_380 = retime_s1_144_reg_reg_N30;
 reg retime_s1_145_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_145_reg_reg_N30 <= n_1435;
 assign n_382 = retime_s1_145_reg_reg_N30;
 reg retime_s1_146_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_146_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_39;
 assign n_384 = retime_s1_146_reg_reg_N30;
 reg retime_s1_147_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_147_reg_reg_N30 <= n_596;
 assign n_386 = retime_s1_147_reg_reg_N30;
 reg retime_s1_148_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s1_148_reg_reg_N30 <= n_595;
 assign n_387 = retime_s1_148_reg_reg_N30;
 reg retime_s1_149_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_149_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_223;
 assign n_389 = retime_s1_149_reg_reg_N30;
 reg retime_s1_150_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_150_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_2;
 assign n_391 = retime_s1_150_reg_reg_N30;
 reg retime_s1_151_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_151_reg_reg_N30 <= n_1433;
 assign n_393 = retime_s1_151_reg_reg_N30;
 reg retime_s1_152_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_152_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_7;
 assign n_395 = retime_s1_152_reg_reg_N30;
 reg retime_s1_153_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_153_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_225;
 assign n_397 = retime_s1_153_reg_reg_N30;
 reg retime_s1_154_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_154_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_225;
 assign n_398 = retime_s1_154_reg_reg_N30;
 reg retime_s1_155_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_155_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_344;
 assign n_399 = retime_s1_155_reg_reg_N30;
 reg retime_s1_156_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_156_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_94;
 assign n_400 = retime_s1_156_reg_reg_N30;
 reg retime_s1_157_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_157_reg_reg_N30 <= csa_tree_add_86_2_n_29;
 assign n_401 = retime_s1_157_reg_reg_N30;
 reg retime_s1_158_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_158_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_44;
 assign n_402 = retime_s1_158_reg_reg_N30;
 reg retime_s1_159_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_159_reg_reg_N30 <= n_1442;
 assign n_403 = retime_s1_159_reg_reg_N30;
 reg retime_s1_160_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_160_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_42;
 assign n_404 = retime_s1_160_reg_reg_N30;
 reg retime_s1_161_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_161_reg_reg_N30 <= csa_tree_add_86_2_n_6;
 assign n_405 = retime_s1_161_reg_reg_N30;
 reg retime_s1_162_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_162_reg_reg_N30 <= {in5[1]};
 assign n_406 = retime_s1_162_reg_reg_N30;
 reg retime_s1_163_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_163_reg_reg_N30 <= n_660;
 assign n_407 = retime_s1_163_reg_reg_N30;
 reg retime_s1_164_reg_reg_N30;
 always @(posedge clk)
         retime_s1_164_reg_reg_N30 <= n_1021;
 assign n_408 = retime_s1_164_reg_reg_N30;
 reg retime_s1_165_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_165_reg_reg_N30 <= csa_tree_add_86_2_n_26;
 assign n_409 = retime_s1_165_reg_reg_N30;
 reg retime_s1_166_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_166_reg_reg_N30 <= n_1438;
 assign n_410 = retime_s1_166_reg_reg_N30;
 reg retime_s1_167_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_167_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_45;
 assign n_412 = retime_s1_167_reg_reg_N30;
 reg retime_s1_168_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_168_reg_reg_N30 <= n_1492;
 assign n_414 = retime_s1_168_reg_reg_N30;
 reg retime_s1_169_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_169_reg_reg_N30 <= n_1437;
 assign n_416 = retime_s1_169_reg_reg_N30;
 reg retime_s1_170_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_170_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_38;
 assign n_418 = retime_s1_170_reg_reg_N30;
 reg retime_s1_171_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_171_reg_reg_N30 <= csa_tree_add_86_2_n_28;
 assign n_420 = retime_s1_171_reg_reg_N30;
 reg retime_s1_172_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_172_reg_reg_N30 <= n_1446;
 assign n_421 = retime_s1_172_reg_reg_N30;
 reg retime_s1_173_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_173_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_40;
 assign n_422 = retime_s1_173_reg_reg_N30;
 reg retime_s1_174_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_174_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_221;
 assign n_423 = retime_s1_174_reg_reg_N30;
 reg retime_s1_175_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_175_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_4;
 assign n_424 = retime_s1_175_reg_reg_N30;
 reg retime_s1_176_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_176_reg_reg_N30 <= {in5[3]};
 assign n_425 = retime_s1_176_reg_reg_N30;
 reg retime_s1_177_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_177_reg_reg_N30 <= csa_tree_add_86_2_n_4;
 assign n_426 = retime_s1_177_reg_reg_N30;
 reg retime_s1_178_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_178_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_343;
 assign n_427 = retime_s1_178_reg_reg_N30;
 reg retime_s1_179_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_179_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_43;
 assign n_428 = retime_s1_179_reg_reg_N30;
 reg retime_s1_180_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_180_reg_reg_N30 <= n_1499;
 assign n_429 = retime_s1_180_reg_reg_N30;
 reg retime_s1_181_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_181_reg_reg_N30 <= {in5[0]};
 assign n_430 = retime_s1_181_reg_reg_N30;
 reg retime_s1_182_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_182_reg_reg_N30 <= csa_tree_add_86_2_n_5;
 assign n_431 = retime_s1_182_reg_reg_N30;
 reg retime_s1_183_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s1_183_reg_reg_N30 <= n_536;
 assign n_432 = retime_s1_183_reg_reg_N30;
 reg retime_s1_184_reg_reg_N30;
 always @(posedge clk)
         retime_s1_184_reg_reg_N30 <= n_790;
 assign csa_tree_add_106_2_groupi_n_337 = retime_s1_184_reg_reg_N30;
 reg retime_s1_185_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_185_reg_reg_N30 <= csa_tree_add_86_2_n_7;
 assign n_434 = retime_s1_185_reg_reg_N30;
 reg retime_s1_186_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_186_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_1;
 assign n_435 = retime_s1_186_reg_reg_N30;
 reg retime_s1_187_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_187_reg_reg_N30 <= n_987;
 assign n_436 = retime_s1_187_reg_reg_N30;
 reg retime_s1_188_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_188_reg_reg_N30 <= n_795;
 assign n_437 = retime_s1_188_reg_reg_N30;
 reg retime_s1_189_reg_reg_N30;
 always @(posedge clk)
         retime_s1_189_reg_reg_N30 <= n_594;
 assign n_438 = retime_s1_189_reg_reg_N30;
 reg retime_s1_190_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_190_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_41;
 assign n_439 = retime_s1_190_reg_reg_N30;
 reg retime_s1_191_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_191_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_226;
 assign n_440 = retime_s1_191_reg_reg_N30;
 reg retime_s1_192_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_192_reg_reg_N30 <= csa_tree_add_106_2_groupi_n_226;
 assign n_441 = retime_s1_192_reg_reg_N30;
 reg retime_s1_193_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_193_reg_reg_N30 <= n_590;
 assign n_442 = retime_s1_193_reg_reg_N30;
 reg retime_s1_194_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s1_194_reg_reg_N30 <= n_654;
 assign n_443 = retime_s1_194_reg_reg_N30;
 reg retime_s1_195_reg_reg_N30;
 always @(posedge clk)
         retime_s1_195_reg_reg_N30 <= n_216;
 assign n_444 = retime_s1_195_reg_reg_N30;
 reg retime_s2_1_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_1_reg_reg_N30 <= n_0;
 assign n_1 = retime_s2_1_reg_reg_N30;
 reg retime_s2_2_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_2_reg_reg_N30 <= n_1380;
 assign n_3 = retime_s2_2_reg_reg_N30;
 reg retime_s2_3_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_3_reg_reg_N30 <= n_1352;
 assign n_4 = retime_s2_3_reg_reg_N30;
 reg retime_s2_4_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_4_reg_reg_N30 <= n_1008;
 assign n_5 = retime_s2_4_reg_reg_N30;
 reg retime_s2_5_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_5_reg_reg_N30 <= n_258;
 assign n_6 = retime_s2_5_reg_reg_N30;
 reg retime_s2_6_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_6_reg_reg_N30 <= n_778;
 assign n_7 = retime_s2_6_reg_reg_N30;
 reg retime_s2_7_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_7_reg_reg_N30 <= n_976;
 assign n_9 = retime_s2_7_reg_reg_N30;
 reg retime_s2_8_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_8_reg_reg_N30 <= n_975;
 assign n_10 = retime_s2_8_reg_reg_N30;
 reg retime_s2_9_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_9_reg_reg_N30 <= n_482;
 assign n_11 = retime_s2_9_reg_reg_N30;
 reg retime_s2_10_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_10_reg_reg_N30 <= n_478;
 assign n_12 = retime_s2_10_reg_reg_N30;
 reg retime_s2_11_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_11_reg_reg_N30 <= n_472;
 assign n_13 = retime_s2_11_reg_reg_N30;
 reg retime_s2_12_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_12_reg_reg_N30 <= n_486;
 assign n_14 = retime_s2_12_reg_reg_N30;
 reg retime_s2_13_reg_reg_N30;
 always @(posedge clk)
         retime_s2_13_reg_reg_N30 <= n_556;
 assign n_15 = retime_s2_13_reg_reg_N30;
 reg retime_s2_14_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_14_reg_reg_N30 <= n_576;
 assign n_16 = retime_s2_14_reg_reg_N30;
 reg retime_s2_15_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s2_15_reg_reg_N30 <= n_699;
 assign n_17 = retime_s2_15_reg_reg_N30;
 reg retime_s2_16_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s2_16_reg_reg_N30 <= n_698;
 assign n_18 = retime_s2_16_reg_reg_N30;
 reg retime_s2_17_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_17_reg_reg_N30 <= n_468;
 assign n_19 = retime_s2_17_reg_reg_N30;
 reg retime_s2_18_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_18_reg_reg_N30 <= n_460;
 assign n_20 = retime_s2_18_reg_reg_N30;
 reg retime_s2_19_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_19_reg_reg_N30 <= n_579;
 assign n_21 = retime_s2_19_reg_reg_N30;
 reg retime_s2_20_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_20_reg_reg_N30 <= n_578;
 assign n_22 = retime_s2_20_reg_reg_N30;
 reg retime_s2_21_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_21_reg_reg_N30 <= n_455;
 assign n_23 = retime_s2_21_reg_reg_N30;
 reg retime_s2_22_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_22_reg_reg_N30 <= n_451;
 assign n_24 = retime_s2_22_reg_reg_N30;
 reg retime_s2_23_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_23_reg_reg_N30 <= n_986;
 assign n_25 = retime_s2_23_reg_reg_N30;
 reg retime_s2_24_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_24_reg_reg_N30 <= n_449;
 assign n_26 = retime_s2_24_reg_reg_N30;
 reg retime_s2_25_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_25_reg_reg_N30 <= n_1007;
 assign n_27 = retime_s2_25_reg_reg_N30;
 reg retime_s2_26_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_26_reg_reg_N30 <= n_1006;
 assign n_28 = retime_s2_26_reg_reg_N30;
 reg retime_s2_27_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_27_reg_reg_N30 <= n_447;
 assign n_29 = retime_s2_27_reg_reg_N30;
 reg retime_s2_28_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_28_reg_reg_N30 <= n_446;
 assign n_30 = retime_s2_28_reg_reg_N30;
 reg retime_s2_29_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_29_reg_reg_N30 <= n_445;
 assign n_31 = retime_s2_29_reg_reg_N30;
 reg retime_s2_30_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_30_reg_reg_N30 <= n_941;
 assign n_32 = retime_s2_30_reg_reg_N30;
 reg retime_s2_31_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_31_reg_reg_N30 <= n_940;
 assign n_33 = retime_s2_31_reg_reg_N30;
 reg retime_s2_32_reg_reg_N30;
 always @(posedge clk)
         retime_s2_32_reg_reg_N30 <= n_457;
 assign mul_109_11_n_41 = retime_s2_32_reg_reg_N30;
 reg retime_s2_33_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_33_reg_reg_N30 <= n_470;
 assign n_34 = retime_s2_33_reg_reg_N30;
 reg retime_s2_34_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_34_reg_reg_N30 <= n_184;
 assign n_35 = retime_s2_34_reg_reg_N30;
 reg retime_s2_35_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_35_reg_reg_N30 <= n_183;
 assign n_36 = retime_s2_35_reg_reg_N30;
 reg retime_s2_36_reg_reg_N30;
 always @(posedge clk)
         retime_s2_36_reg_reg_N30 <= n_464;
 assign mul_109_11_n_25 = retime_s2_36_reg_reg_N30;
 reg retime_s2_37_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_37_reg_reg_N30 <= n_462;
 assign n_37 = retime_s2_37_reg_reg_N30;
 reg retime_s2_38_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_38_reg_reg_N30 <= n_182;
 assign n_38 = retime_s2_38_reg_reg_N30;
 reg retime_s2_39_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_39_reg_reg_N30 <= n_181;
 assign n_39 = retime_s2_39_reg_reg_N30;
 reg retime_s2_40_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_40_reg_reg_N30 <= n_1013;
 assign n_40 = retime_s2_40_reg_reg_N30;
 reg retime_s2_41_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_41_reg_reg_N30 <= n_668;
 assign n_41 = retime_s2_41_reg_reg_N30;
 reg retime_s2_42_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_42_reg_reg_N30 <= n_186;
 assign n_42 = retime_s2_42_reg_reg_N30;
 reg retime_s2_43_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_43_reg_reg_N30 <= n_185;
 assign n_43 = retime_s2_43_reg_reg_N30;
 reg retime_s2_44_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_44_reg_reg_N30 <= n_454;
 assign n_44 = retime_s2_44_reg_reg_N30;
 reg retime_s2_45_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_45_reg_reg_N30 <= n_453;
 assign n_45 = retime_s2_45_reg_reg_N30;
 reg retime_s2_46_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_46_reg_reg_N30 <= n_188;
 assign n_46 = retime_s2_46_reg_reg_N30;
 reg retime_s2_47_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_47_reg_reg_N30 <= n_694;
 assign n_47 = retime_s2_47_reg_reg_N30;
 reg retime_s2_48_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_48_reg_reg_N30 <= n_581;
 assign n_48 = retime_s2_48_reg_reg_N30;
 reg retime_s2_49_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_49_reg_reg_N30 <= n_539;
 assign n_49 = retime_s2_49_reg_reg_N30;
 reg retime_s2_50_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s2_50_reg_reg_N30 <= n_538;
 assign n_50 = retime_s2_50_reg_reg_N30;
 reg retime_s2_51_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_51_reg_reg_N30 <= n_978;
 assign n_51 = retime_s2_51_reg_reg_N30;
 reg retime_s2_52_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_52_reg_reg_N30 <= n_977;
 assign n_52 = retime_s2_52_reg_reg_N30;
 reg retime_s2_53_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s2_53_reg_reg_N30 <= n_192;
 assign n_53 = retime_s2_53_reg_reg_N30;
 reg retime_s2_54_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s2_54_reg_reg_N30 <= n_191;
 assign n_54 = retime_s2_54_reg_reg_N30;
 reg retime_s2_55_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_55_reg_reg_N30 <= n_189;
 assign n_55 = retime_s2_55_reg_reg_N30;
 reg retime_s2_56_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s2_56_reg_reg_N30 <= n_672;
 assign n_56 = retime_s2_56_reg_reg_N30;
 reg retime_s2_57_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s2_57_reg_reg_N30 <= n_671;
 assign n_57 = retime_s2_57_reg_reg_N30;
 reg retime_s2_58_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s2_58_reg_reg_N30 <= n_194;
 assign n_58 = retime_s2_58_reg_reg_N30;
 reg retime_s2_59_reg_reg_N30;
 always @(posedge clk)
         if (n_465)
         retime_s2_59_reg_reg_N30 <= n_193;
 assign n_59 = retime_s2_59_reg_reg_N30;
 reg retime_s2_60_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_60_reg_reg_N30 <= n_474;
 assign n_60 = retime_s2_60_reg_reg_N30;
 reg retime_s2_61_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_61_reg_reg_N30 <= n_476;
 assign n_61 = retime_s2_61_reg_reg_N30;
 reg retime_s2_62_reg_reg_N30;
 always @(posedge clk)
         retime_s2_62_reg_reg_N30 <= n_573;
 assign n_62 = retime_s2_62_reg_reg_N30;
 reg retime_s2_63_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_63_reg_reg_N30 <= n_1050;
 assign n_63 = retime_s2_63_reg_reg_N30;
 reg retime_s2_64_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_64_reg_reg_N30 <= n_1051;
 assign n_64 = retime_s2_64_reg_reg_N30;
 reg retime_s2_65_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_65_reg_reg_N30 <= n_1060;
 assign n_65 = retime_s2_65_reg_reg_N30;
 reg retime_s2_66_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_66_reg_reg_N30 <= n_1053;
 assign n_66 = retime_s2_66_reg_reg_N30;
 reg retime_s2_67_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_67_reg_reg_N30 <= n_717;
 assign n_67 = retime_s2_67_reg_reg_N30;
 reg retime_s2_68_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_68_reg_reg_N30 <= n_683;
 assign n_68 = retime_s2_68_reg_reg_N30;
 reg retime_s2_69_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_69_reg_reg_N30 <= n_673;
 assign n_69 = retime_s2_69_reg_reg_N30;
 reg retime_s2_70_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_70_reg_reg_N30 <= n_973;
 assign n_70 = retime_s2_70_reg_reg_N30;
 reg retime_s2_71_reg_reg_N30;
 always @(posedge clk)
         retime_s2_71_reg_reg_N30 <= n_708;
 assign n_71 = retime_s2_71_reg_reg_N30;
 reg retime_s2_72_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_72_reg_reg_N30 <= n_1042;
 assign n_72 = retime_s2_72_reg_reg_N30;
 reg retime_s2_73_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_73_reg_reg_N30 <= n_497;
 assign n_73 = retime_s2_73_reg_reg_N30;
 reg retime_s2_74_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_74_reg_reg_N30 <= n_490;
 assign n_74 = retime_s2_74_reg_reg_N30;
 reg retime_s2_75_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_75_reg_reg_N30 <= n_504;
 assign n_75 = retime_s2_75_reg_reg_N30;
 reg retime_s2_76_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_76_reg_reg_N30 <= n_717;
 assign n_76 = retime_s2_76_reg_reg_N30;
 reg retime_s2_77_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_77_reg_reg_N30 <= n_480;
 assign n_77 = retime_s2_77_reg_reg_N30;
 reg retime_s2_78_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_78_reg_reg_N30 <= n_484;
 assign n_79 = retime_s2_78_reg_reg_N30;
 reg retime_s2_79_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_79_reg_reg_N30 <= n_1010;
 assign n_80 = retime_s2_79_reg_reg_N30;
 reg retime_s2_80_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_80_reg_reg_N30 <= n_488;
 assign n_81 = retime_s2_80_reg_reg_N30;
 reg retime_s2_81_reg_reg_N30;
 always @(posedge clk)
         retime_s2_81_reg_reg_N30 <= n_494;
 assign mul_109_11_n_39 = retime_s2_81_reg_reg_N30;
 reg retime_s2_82_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_82_reg_reg_N30 <= n_503;
 assign n_82 = retime_s2_82_reg_reg_N30;
 reg retime_s2_83_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_83_reg_reg_N30 <= n_500;
 assign n_83 = retime_s2_83_reg_reg_N30;
 reg retime_s2_84_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_84_reg_reg_N30 <= n_492;
 assign n_84 = retime_s2_84_reg_reg_N30;
 reg retime_s2_85_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_85_reg_reg_N30 <= n_949;
 assign n_85 = retime_s2_85_reg_reg_N30;
 reg retime_s2_86_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_86_reg_reg_N30 <= n_499;
 assign n_86 = retime_s2_86_reg_reg_N30;
 reg retime_s2_87_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_87_reg_reg_N30 <= n_514;
 assign n_87 = retime_s2_87_reg_reg_N30;
 reg retime_s2_88_reg_reg_N30;
 always @(posedge clk)
         retime_s2_88_reg_reg_N30 <= n_508;
 assign mul_109_11_n_393 = retime_s2_88_reg_reg_N30;
 reg retime_s2_89_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_89_reg_reg_N30 <= n_520;
 assign n_88 = retime_s2_89_reg_reg_N30;
 reg retime_s2_90_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_90_reg_reg_N30 <= n_89;
 assign n_90 = retime_s2_90_reg_reg_N30;
 reg retime_s2_91_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_91_reg_reg_N30 <= n_1158;
 assign n_92 = retime_s2_91_reg_reg_N30;
 reg retime_s2_92_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_92_reg_reg_N30 <= n_1157;
 assign n_95 = retime_s2_92_reg_reg_N30;
 reg retime_s2_93_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_93_reg_reg_N30 <= n_958;
 assign n_96 = retime_s2_93_reg_reg_N30;
 reg retime_s2_94_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_94_reg_reg_N30 <= n_658;
 assign n_97 = retime_s2_94_reg_reg_N30;
 reg retime_s2_95_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_95_reg_reg_N30 <= n_558;
 assign n_98 = retime_s2_95_reg_reg_N30;
 reg retime_s2_96_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_96_reg_reg_N30 <= n_532;
 assign n_99 = retime_s2_96_reg_reg_N30;
 reg retime_s2_97_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_97_reg_reg_N30 <= n_521;
 assign n_100 = retime_s2_97_reg_reg_N30;
 reg retime_s2_98_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_98_reg_reg_N30 <= n_511;
 assign n_101 = retime_s2_98_reg_reg_N30;
 reg retime_s2_99_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_99_reg_reg_N30 <= n_245;
 assign n_102 = retime_s2_99_reg_reg_N30;
 reg retime_s2_100_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_100_reg_reg_N30 <= n_105;
 assign n_106 = retime_s2_100_reg_reg_N30;
 reg retime_s2_101_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_101_reg_reg_N30 <= n_552;
 assign n_135 = retime_s2_101_reg_reg_N30;
 reg retime_s2_102_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_102_reg_reg_N30 <= n_604;
 assign n_136 = retime_s2_102_reg_reg_N30;
 reg retime_s2_103_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_103_reg_reg_N30 <= n_171;
 assign n_310 = retime_s2_103_reg_reg_N30;
 reg retime_s2_104_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_104_reg_reg_N30 <= n_246;
 assign n_311 = retime_s2_104_reg_reg_N30;
 reg retime_s2_105_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_105_reg_reg_N30 <= n_361;
 assign n_362 = retime_s2_105_reg_reg_N30;
 reg retime_s2_106_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_106_reg_reg_N30 <= n_369;
 assign n_370 = retime_s2_106_reg_reg_N30;
 reg retime_s2_107_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_107_reg_reg_N30 <= n_378;
 assign n_379 = retime_s2_107_reg_reg_N30;
 reg retime_s2_108_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_108_reg_reg_N30 <= n_380;
 assign n_381 = retime_s2_108_reg_reg_N30;
 reg retime_s2_109_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_109_reg_reg_N30 <= n_382;
 assign n_383 = retime_s2_109_reg_reg_N30;
 reg retime_s2_110_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_110_reg_reg_N30 <= n_384;
 assign n_385 = retime_s2_110_reg_reg_N30;
 reg retime_s2_111_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_111_reg_reg_N30 <= n_387;
 assign n_388 = retime_s2_111_reg_reg_N30;
 reg retime_s2_112_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_112_reg_reg_N30 <= n_389;
 assign n_390 = retime_s2_112_reg_reg_N30;
 reg retime_s2_113_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_113_reg_reg_N30 <= n_391;
 assign n_392 = retime_s2_113_reg_reg_N30;
 reg retime_s2_114_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_114_reg_reg_N30 <= n_393;
 assign n_394 = retime_s2_114_reg_reg_N30;
 reg retime_s2_115_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_115_reg_reg_N30 <= n_395;
 assign n_396 = retime_s2_115_reg_reg_N30;
 reg retime_s2_116_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_116_reg_reg_N30 <= n_410;
 assign n_411 = retime_s2_116_reg_reg_N30;
 reg retime_s2_117_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_117_reg_reg_N30 <= n_412;
 assign n_413 = retime_s2_117_reg_reg_N30;
 reg retime_s2_118_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_118_reg_reg_N30 <= n_414;
 assign n_415 = retime_s2_118_reg_reg_N30;
 reg retime_s2_119_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_119_reg_reg_N30 <= n_416;
 assign n_417 = retime_s2_119_reg_reg_N30;
 reg retime_s2_120_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_120_reg_reg_N30 <= n_418;
 assign n_419 = retime_s2_120_reg_reg_N30;
 reg retime_s2_121_reg_reg_N30;
 always @(posedge clk)
         if (stall == 1'B0)
         retime_s2_121_reg_reg_N30 <= n_432;
 assign n_433 = retime_s2_121_reg_reg_N30;
 assign add_57_2_n_2 = ~(add_57_2_n_21 & (add_57_2_n_26 & ~add_57_2_n_38));
 assign n_1315 = (add_57_2_n_48 ^ add_57_2_n_16);
 assign add_57_2_n_48 = ~(add_57_2_n_44 | ~add_57_2_n_12);
 assign n_1314 = ~(add_57_2_n_2 & (add_57_2_n_7 & add_57_2_n_31));
 assign n_1316 = ~(add_57_2_n_42 ^ add_57_2_n_18);
 assign n_1317 = ~(add_57_2_n_43 ^ add_57_2_n_17);
 assign add_57_2_n_44 = ~(add_57_2_n_42 | add_57_2_n_3);
 assign add_57_2_n_43 = ~(add_57_2_n_40 | ~add_57_2_n_11);
 assign add_57_2_n_42 = ~(add_57_2_n_39 | add_57_2_n_27);
 assign n_1318 = ~(add_57_2_n_38 ^ add_57_2_n_23);
 assign add_57_2_n_40 = ~(add_57_2_n_38 | add_57_2_n_13);
 assign add_57_2_n_39 = ~(add_57_2_n_38 | ~add_57_2_n_21);
 assign add_57_2_n_38 = ~(add_57_2_n_36 | add_57_2_n_8);
 assign n_1319 = ~(add_57_2_n_34 ^ add_57_2_n_24);
 assign add_57_2_n_36 = ~(add_57_2_n_35 | add_57_2_n_15);
 assign add_57_2_n_35 = ~(add_57_2_n_32 | add_57_2_n_0);
 assign add_57_2_n_34 = ~(add_57_2_n_0 | ~(add_57_2_n_30 | add_57_2_n_4));
 assign n_1320 = ~(add_57_2_n_30 ^ add_57_2_n_19);
 assign add_57_2_n_32 = ~(add_57_2_n_30 | add_57_2_n_4);
 assign add_57_2_n_31 = ~(add_57_2_n_25 | (add_57_2_n_27 & add_57_2_n_26));
 assign add_57_2_n_30 = ~(add_57_2_n_28 | add_57_2_n_1);
 assign n_1321 = (add_57_2_n_22 ^ add_57_2_n_6);
 assign add_57_2_n_28 = ~(add_57_2_n_9 | add_57_2_n_6);
 assign add_57_2_n_27 = ~(add_57_2_n_10 & (add_57_2_n_5 | add_57_2_n_11));
 assign add_57_2_n_25 = ~(add_57_2_n_14 | add_57_2_n_12);
 assign add_57_2_n_24 = ~(add_57_2_n_15 | add_57_2_n_8);
 assign add_57_2_n_23 = ~(add_57_2_n_13 | ~add_57_2_n_11);
 assign add_57_2_n_22 = (add_57_2_n_9 | add_57_2_n_1);
 assign add_57_2_n_26 = ~(add_57_2_n_3 | add_57_2_n_14);
 assign n_1322 = ({in8[0]} ^ {in7[0]});
 assign add_57_2_n_21 = ~(add_57_2_n_13 | add_57_2_n_5);
 assign add_57_2_n_19 = ~(add_57_2_n_4 | add_57_2_n_0);
 assign add_57_2_n_18 = ~(add_57_2_n_3 | ~add_57_2_n_12);
 assign add_57_2_n_17 = ~(add_57_2_n_5 | ~add_57_2_n_10);
 assign add_57_2_n_16 = ~(add_57_2_n_7 & ~add_57_2_n_14);
 assign add_57_2_n_15 = ~({in8[3]} | {in7[3]});
 assign add_57_2_n_14 = ~({in8[7]} | {in7[7]});
 assign add_57_2_n_13 = ~({in8[4]} | {in7[4]});
 assign add_57_2_n_12 = ~({in8[6]} & {in7[6]});
 assign add_57_2_n_11 = ~({in8[4]} & {in7[4]});
 assign add_57_2_n_10 = ~({in8[5]} & {in7[5]});
 assign add_57_2_n_9 = ~({in8[1]} | {in7[1]});
 assign add_57_2_n_8 = ({in8[3]} & {in7[3]});
 assign add_57_2_n_7 = ~({in8[7]} & {in7[7]});
 assign add_57_2_n_6 = ~({in8[0]} & {in7[0]});
 assign add_57_2_n_5 = ~({in8[5]} | {in7[5]});
 assign add_57_2_n_4 = ~({in8[2]} | {in7[2]});
 assign add_57_2_n_3 = ~({in8[6]} | {in7[6]});
 assign add_57_2_n_1 = ({in8[1]} & {in7[1]});
 assign add_57_2_n_0 = ({in8[2]} & {in7[2]});
 assign add_100_2_n_40 = ~(add_100_2_n_8 & (add_100_2_n_34 | add_100_2_n_0));
 assign n_1439 = ~(add_100_2_n_24 & (add_100_2_n_36 & (add_100_2_n_6 | add_100_2_n_8)));
 assign n_1441 = ~(add_100_2_n_34 ^ add_100_2_n_14);
 assign add_100_2_n_36 = ~(add_100_2_n_5 | (add_100_2_n_32 & (add_100_2_n_16 & add_100_2_n_18)));
 assign add_100_2_n_35 = ~(add_100_2_n_11 & (add_100_2_n_31 | add_100_2_n_7));
 assign add_100_2_n_34 = ~(add_100_2_n_21 | (add_100_2_n_32 & add_100_2_n_16));
 assign n_1443 = ~(add_100_2_n_31 ^ add_100_2_n_20);
 assign add_100_2_n_31 = ~add_100_2_n_32;
 assign add_100_2_n_32 = ~(add_100_2_n_4 & (add_100_2_n_29 | add_100_2_n_12));
 assign add_100_2_n_29 = ~(add_100_2_n_9 | (add_100_2_n_26 & add_100_2_n_2));
 assign add_100_2_n_28 = ~(add_100_2_n_10 & ~(add_100_2_n_26 & add_100_2_n_2));
 assign n_1445 = ~(add_100_2_n_26 ^ add_100_2_n_15);
 assign add_100_2_n_24 = ~(add_100_2_n_21 & add_100_2_n_18);
 assign add_100_2_n_22 = ({in4[0]} & {in3[0]});
 assign n_1447 = ({in4[0]} ^ {in3[0]});
 assign add_100_2_n_21 = ~(add_100_2_n_3 & (add_100_2_n_1 | add_100_2_n_11));
 assign add_100_2_n_20 = ~(add_100_2_n_7 | ~add_100_2_n_11);
 assign add_100_2_n_19 = ~(add_100_2_n_4 & ~add_100_2_n_12);
 assign add_100_2_n_18 = ~(add_100_2_n_0 | add_100_2_n_6);
 assign add_100_2_n_17 = (add_100_2_n_6 | add_100_2_n_5);
 assign add_100_2_n_16 = ~(add_100_2_n_7 | add_100_2_n_1);
 assign add_100_2_n_15 = ~(add_100_2_n_2 & add_100_2_n_10);
 assign add_100_2_n_14 = ~(add_100_2_n_0 | ~add_100_2_n_8);
 assign add_100_2_n_13 = ~(add_100_2_n_3 & ~add_100_2_n_1);
 assign add_100_2_n_9 = ~add_100_2_n_10;
 assign add_100_2_n_12 = ~({in4[3]} | {in3[3]});
 assign add_100_2_n_11 = ~({in4[4]} & {in3[4]});
 assign add_100_2_n_10 = ~({in4[2]} & {in3[2]});
 assign add_100_2_n_8 = ~({in4[6]} & {in3[6]});
 assign add_100_2_n_7 = ~({in4[4]} | {in3[4]});
 assign add_100_2_n_6 = ~({in4[7]} | {in3[7]});
 assign add_100_2_n_5 = ({in4[7]} & {in3[7]});
 assign add_100_2_n_4 = ~({in4[3]} & {in3[3]});
 assign add_100_2_n_3 = ~({in4[5]} & {in3[5]});
 assign add_100_2_n_2 = ({in4[2]} | {in3[2]});
 assign add_100_2_n_1 = ~({in4[5]} | {in3[5]});
 assign add_100_2_n_0 = ~({in4[6]} | {in3[6]});
 assign csa_tree_add_64_2_groupi_n_11 = (csa_tree_add_64_2_groupi_n_12 | csa_tree_add_64_2_groupi_n_61);
 assign n_1274 = (csa_tree_add_64_2_groupi_n_72 & csa_tree_add_64_2_groupi_n_28);
 assign n_1275 = (csa_tree_add_64_2_groupi_n_72 ^ csa_tree_add_64_2_groupi_n_28);
 assign n_1276 = ~(csa_tree_add_64_2_groupi_n_83 & ~csa_tree_add_64_2_groupi_n_82);
 assign csa_tree_add_64_2_groupi_n_83 = ~(csa_tree_add_64_2_groupi_n_81 & csa_tree_add_64_2_groupi_n_59);
 assign csa_tree_add_64_2_groupi_n_82 = ~(csa_tree_add_64_2_groupi_n_78 | (csa_tree_add_64_2_groupi_n_43
    | csa_tree_add_64_2_groupi_n_59));
 assign csa_tree_add_64_2_groupi_n_81 = ~(csa_tree_add_64_2_groupi_n_77 & csa_tree_add_64_2_groupi_n_42);
 assign n_1277 = ~(csa_tree_add_64_2_groupi_n_76 & ~csa_tree_add_64_2_groupi_n_75);
 assign n_1278 = ~(csa_tree_add_64_2_groupi_n_74 & ~csa_tree_add_64_2_groupi_n_73);
 assign csa_tree_add_64_2_groupi_n_78 = ~csa_tree_add_64_2_groupi_n_77;
 assign csa_tree_add_64_2_groupi_n_77 = ~(csa_tree_add_64_2_groupi_n_47 & (csa_tree_add_64_2_groupi_n_12
    | csa_tree_add_64_2_groupi_n_61));
 assign csa_tree_add_64_2_groupi_n_76 = ~(csa_tree_add_64_2_groupi_n_11 & csa_tree_add_64_2_groupi_n_58);
 assign csa_tree_add_64_2_groupi_n_75 = ~(csa_tree_add_64_2_groupi_n_12 | (csa_tree_add_64_2_groupi_n_61
    | csa_tree_add_64_2_groupi_n_58));
 assign csa_tree_add_64_2_groupi_n_74 = ~(csa_tree_add_64_2_groupi_n_10 & csa_tree_add_64_2_groupi_n_57);
 assign csa_tree_add_64_2_groupi_n_73 = ~(csa_tree_add_64_2_groupi_n_5 | (csa_tree_add_64_2_groupi_n_40
    | csa_tree_add_64_2_groupi_n_57));
 assign csa_tree_add_64_2_groupi_n_72 = ~(csa_tree_add_64_2_groupi_n_67 & (csa_tree_add_64_2_groupi_n_71
    | (csa_tree_add_64_2_groupi_n_6 | csa_tree_add_64_2_groupi_n_55)));
 assign csa_tree_add_64_2_groupi_n_71 = ~(csa_tree_add_64_2_groupi_n_69 | csa_tree_add_64_2_groupi_n_3);
 assign n_1280 = ~(csa_tree_add_64_2_groupi_n_13 ^ csa_tree_add_64_2_groupi_n_62);
 assign csa_tree_add_64_2_groupi_n_69 = ~(csa_tree_add_64_2_groupi_n_13 | csa_tree_add_64_2_groupi_n_53);
 assign csa_tree_add_64_2_groupi_n_67 = ~(csa_tree_add_64_2_groupi_n_60 | (csa_tree_add_64_2_groupi_n_61
    & csa_tree_add_64_2_groupi_n_54));
 assign csa_tree_add_64_2_groupi_n_64 = ((csa_tree_add_64_2_groupi_n_34 & n_1480) | ((n_1480 & {in4[1]})
    | ({in4[1]} & csa_tree_add_64_2_groupi_n_34)));
 assign n_1282 = (n_1480 ^ ({in4[1]} ^ csa_tree_add_64_2_groupi_n_34));
 assign csa_tree_add_64_2_groupi_n_62 = ~((csa_tree_add_64_2_groupi_n_14 & ~csa_tree_add_64_2_groupi_n_31)
    | (csa_tree_add_64_2_groupi_n_50 & csa_tree_add_64_2_groupi_n_31));
 assign csa_tree_add_64_2_groupi_n_61 = ~(csa_tree_add_64_2_groupi_n_45 & (csa_tree_add_64_2_groupi_n_49
    | csa_tree_add_64_2_groupi_n_41));
 assign csa_tree_add_64_2_groupi_n_60 = ~(csa_tree_add_64_2_groupi_n_44 & (csa_tree_add_64_2_groupi_n_48
    | csa_tree_add_64_2_groupi_n_42));
 assign csa_tree_add_64_2_groupi_n_59 = ~(csa_tree_add_64_2_groupi_n_44 & ~csa_tree_add_64_2_groupi_n_48);
 assign csa_tree_add_64_2_groupi_n_58 = ~(csa_tree_add_64_2_groupi_n_42 & ~csa_tree_add_64_2_groupi_n_46);
 assign csa_tree_add_64_2_groupi_n_57 = ~(csa_tree_add_64_2_groupi_n_45 & ~csa_tree_add_64_2_groupi_n_49);
 assign csa_tree_add_64_2_groupi_n_56 = ~(csa_tree_add_64_2_groupi_n_40 | ~csa_tree_add_64_2_groupi_n_4);
 assign csa_tree_add_64_2_groupi_n_55 = ~csa_tree_add_64_2_groupi_n_54;
 assign csa_tree_add_64_2_groupi_n_54 = ~(csa_tree_add_64_2_groupi_n_46 | csa_tree_add_64_2_groupi_n_48);
 assign csa_tree_add_64_2_groupi_n_53 = ~(csa_tree_add_64_2_groupi_n_31 | csa_tree_add_64_2_groupi_n_50);
 assign csa_tree_add_64_2_groupi_n_52 = ~csa_tree_add_64_2_groupi_n_51;
 assign csa_tree_add_64_2_groupi_n_51 = ~(csa_tree_add_64_2_groupi_n_27 | csa_tree_add_64_2_groupi_n_2);
 assign csa_tree_add_64_2_groupi_n_50 = ~csa_tree_add_64_2_groupi_n_14;
 assign csa_tree_add_64_2_groupi_n_49 = ~(csa_tree_add_64_2_groupi_n_33 | csa_tree_add_64_2_groupi_n_36);
 assign csa_tree_add_64_2_groupi_n_48 = ~(csa_tree_add_64_2_groupi_n_29 | csa_tree_add_64_2_groupi_n_38);
 assign csa_tree_add_64_2_groupi_n_47 = ~csa_tree_add_64_2_groupi_n_46;
 assign csa_tree_add_64_2_groupi_n_46 = ~(csa_tree_add_64_2_groupi_n_39 | csa_tree_add_64_2_groupi_n_32);
 assign csa_tree_add_64_2_groupi_n_45 = ~(csa_tree_add_64_2_groupi_n_33 & csa_tree_add_64_2_groupi_n_36);
 assign csa_tree_add_64_2_groupi_n_44 = ~(csa_tree_add_64_2_groupi_n_29 & csa_tree_add_64_2_groupi_n_38);
 assign csa_tree_add_64_2_groupi_n_43 = ~csa_tree_add_64_2_groupi_n_42;
 assign csa_tree_add_64_2_groupi_n_42 = ~(csa_tree_add_64_2_groupi_n_39 & csa_tree_add_64_2_groupi_n_32);
 assign csa_tree_add_64_2_groupi_n_40 = ~csa_tree_add_64_2_groupi_n_41;
 assign csa_tree_add_64_2_groupi_n_41 = ~(csa_tree_add_64_2_groupi_n_37 & csa_tree_add_64_2_groupi_n_30);
 assign csa_tree_add_64_2_groupi_n_38 = (({in4[6]} & {in6[6]}) | (({in6[6]} & {in5[6]}) | ({in5[6]} &
    {in4[6]})));
 assign csa_tree_add_64_2_groupi_n_39 = ({in6[6]} ^ ({in5[6]} ^ {in4[6]}));
 assign csa_tree_add_64_2_groupi_n_36 = (({in4[4]} & {in6[4]}) | (({in6[4]} & {in5[4]}) | ({in5[4]} &
    {in4[4]})));
 assign csa_tree_add_64_2_groupi_n_37 = ({in6[4]} ^ ({in5[4]} ^ {in4[4]}));
 assign csa_tree_add_64_2_groupi_n_34 = (({in5[0]} & {in6[0]}) | (({in6[0]} & {in4[0]}) | ({in4[0]} &
    {in5[0]})));
 assign n_1283 = ({in6[0]} ^ ({in4[0]} ^ {in5[0]}));
 assign csa_tree_add_64_2_groupi_n_32 = (({in4[5]} & {in6[5]}) | (({in6[5]} & {in5[5]}) | ({in5[5]} &
    {in4[5]})));
 assign csa_tree_add_64_2_groupi_n_33 = ({in6[5]} ^ ({in5[5]} ^ {in4[5]}));
 assign csa_tree_add_64_2_groupi_n_30 = (({in6[3]} & {in4[3]}) | (({in4[3]} & {in5[3]}) | ({in5[3]} &
    {in6[3]})));
 assign csa_tree_add_64_2_groupi_n_31 = ({in4[3]} ^ ({in5[3]} ^ {in6[3]}));
 assign csa_tree_add_64_2_groupi_n_28 = (({in4[7]} & {in6[7]}) | (({in6[7]} & {in5[7]}) | ({in5[7]} &
    {in4[7]})));
 assign csa_tree_add_64_2_groupi_n_29 = ({in6[7]} ^ ({in5[7]} ^ {in4[7]}));
 assign csa_tree_add_64_2_groupi_n_14 = ~(csa_tree_add_64_2_groupi_n_24 | csa_tree_add_64_2_groupi_n_18);
 assign csa_tree_add_64_2_groupi_n_27 = ~(csa_tree_add_64_2_groupi_n_25 & csa_tree_add_64_2_groupi_n_26);
 assign csa_tree_add_64_2_groupi_n_26 = ~(csa_tree_add_64_2_groupi_n_23 & csa_tree_add_64_2_groupi_n_17);
 assign csa_tree_add_64_2_groupi_n_25 = ~(csa_tree_add_64_2_groupi_n_19 & (csa_tree_add_64_2_groupi_n_20
    & {in5[2]}));
 assign csa_tree_add_64_2_groupi_n_24 = ~(csa_tree_add_64_2_groupi_n_21 | csa_tree_add_64_2_groupi_n_17);
 assign csa_tree_add_64_2_groupi_n_23 = ~(csa_tree_add_64_2_groupi_n_19 & csa_tree_add_64_2_groupi_n_20);
 assign csa_tree_add_64_2_groupi_n_21 = ~({in4[2]} | {in6[2]});
 assign csa_tree_add_64_2_groupi_n_20 = ~(csa_tree_add_64_2_groupi_n_16 & {in4[2]});
 assign csa_tree_add_64_2_groupi_n_19 = ~(csa_tree_add_64_2_groupi_n_15 & {in6[2]});
 assign csa_tree_add_64_2_groupi_n_18 = ~(csa_tree_add_64_2_groupi_n_15 | csa_tree_add_64_2_groupi_n_16);
 assign csa_tree_add_64_2_groupi_n_17 = ~{in5[2]};
 assign csa_tree_add_64_2_groupi_n_16 = ~{in6[2]};
 assign csa_tree_add_64_2_groupi_n_15 = ~{in4[2]};
 assign csa_tree_add_64_2_groupi_n_13 = ~(csa_tree_add_64_2_groupi_n_7 | (csa_tree_add_64_2_groupi_n_64
    & csa_tree_add_64_2_groupi_n_52));
 assign csa_tree_add_64_2_groupi_n_12 = ~(csa_tree_add_64_2_groupi_n_71 | csa_tree_add_64_2_groupi_n_6);
 assign csa_tree_add_64_2_groupi_n_10 = ~(csa_tree_add_64_2_groupi_n_41 & ~csa_tree_add_64_2_groupi_n_5);
 assign n_1279 = ~(csa_tree_add_64_2_groupi_n_71 ^ csa_tree_add_64_2_groupi_n_56);
 assign csa_tree_add_64_2_groupi_n_8 = (csa_tree_add_64_2_groupi_n_7 | csa_tree_add_64_2_groupi_n_51);
 assign csa_tree_add_64_2_groupi_n_7 = (csa_tree_add_64_2_groupi_n_27 & csa_tree_add_64_2_groupi_n_2);
 assign csa_tree_add_64_2_groupi_n_6 = ~(csa_tree_add_64_2_groupi_n_4 & ~csa_tree_add_64_2_groupi_n_49);
 assign csa_tree_add_64_2_groupi_n_5 = ~(csa_tree_add_64_2_groupi_n_71 | ~csa_tree_add_64_2_groupi_n_4);
 assign csa_tree_add_64_2_groupi_n_4 = (csa_tree_add_64_2_groupi_n_37 | csa_tree_add_64_2_groupi_n_30);
 assign csa_tree_add_64_2_groupi_n_3 = ~(csa_tree_add_64_2_groupi_n_14 | ~csa_tree_add_64_2_groupi_n_31);
 assign csa_tree_add_64_2_groupi_n_2 = ({in5[1]} & {in6[1]});
 assign csa_tree_add_71_2_groupi_n_57 = ~csa_tree_add_71_2_groupi_n_108;
 assign csa_tree_add_71_2_groupi_n_56 = csa_tree_add_71_2_groupi_n_4;
 assign n_1284 = (csa_tree_add_71_2_groupi_n_121 & csa_tree_add_71_2_groupi_n_14);
 assign n_1285 = (csa_tree_add_71_2_groupi_n_121 ^ csa_tree_add_71_2_groupi_n_14);
 assign n_1287 = ~(csa_tree_add_71_2_groupi_n_126 & ~csa_tree_add_71_2_groupi_n_125);
 assign n_1286 = ~csa_tree_add_71_2_groupi_n_127;
 assign csa_tree_add_71_2_groupi_n_127 = ~(csa_tree_add_71_2_groupi_n_122 | (csa_tree_add_71_2_groupi_n_111
    & (csa_tree_add_71_2_groupi_n_99 & csa_tree_add_71_2_groupi_n_53)));
 assign csa_tree_add_71_2_groupi_n_126 = ~(csa_tree_add_71_2_groupi_n_120 & csa_tree_add_71_2_groupi_n_88);
 assign csa_tree_add_71_2_groupi_n_125 = ~(csa_tree_add_71_2_groupi_n_117 | (csa_tree_add_71_2_groupi_n_91
    | csa_tree_add_71_2_groupi_n_88));
 assign csa_tree_add_71_2_groupi_n_122 = ~(csa_tree_add_71_2_groupi_n_118 | csa_tree_add_71_2_groupi_n_53);
 assign csa_tree_add_71_2_groupi_n_121 = ~(csa_tree_add_71_2_groupi_n_95 & (csa_tree_add_71_2_groupi_n_108
    | csa_tree_add_71_2_groupi_n_93));
 assign csa_tree_add_71_2_groupi_n_120 = ~(csa_tree_add_71_2_groupi_n_92 & (csa_tree_add_71_2_groupi_n_108
    | csa_tree_add_71_2_groupi_n_81));
 assign csa_tree_add_71_2_groupi_n_119 = ~(csa_tree_add_71_2_groupi_n_62 & (csa_tree_add_71_2_groupi_n_108
    | csa_tree_add_71_2_groupi_n_73));
 assign csa_tree_add_71_2_groupi_n_118 = ~(csa_tree_add_71_2_groupi_n_110 | csa_tree_add_71_2_groupi_n_98);
 assign csa_tree_add_71_2_groupi_n_117 = ~(csa_tree_add_71_2_groupi_n_108 | csa_tree_add_71_2_groupi_n_81);
 assign csa_tree_add_71_2_groupi_n_116 = ~(csa_tree_add_71_2_groupi_n_108 | csa_tree_add_71_2_groupi_n_73);
 assign csa_tree_add_71_2_groupi_n_111 = ~csa_tree_add_71_2_groupi_n_110;
 assign csa_tree_add_71_2_groupi_n_110 = ~(csa_tree_add_71_2_groupi_n_108 | csa_tree_add_71_2_groupi_n_94);
 assign csa_tree_add_71_2_groupi_n_109 = ~(csa_tree_add_71_2_groupi_n_64 & (csa_tree_add_71_2_groupi_n_71
    | csa_tree_add_71_2_groupi_n_103));
 assign csa_tree_add_71_2_groupi_n_108 = ~(csa_tree_add_71_2_groupi_n_89 | csa_tree_add_71_2_groupi_n_105);
 assign csa_tree_add_71_2_groupi_n_105 = ~(csa_tree_add_71_2_groupi_n_71 | (csa_tree_add_71_2_groupi_n_69
    | csa_tree_add_71_2_groupi_n_103));
 assign csa_tree_add_71_2_groupi_n_103 = ~(csa_tree_add_71_2_groupi_n_102 | csa_tree_add_71_2_groupi_n_76);
 assign n_1292 = ~(csa_tree_add_71_2_groupi_n_100 & csa_tree_add_71_2_groupi_n_101);
 assign csa_tree_add_71_2_groupi_n_102 = ~(csa_tree_add_71_2_groupi_n_74 | ~csa_tree_add_71_2_groupi_n_96);
 assign csa_tree_add_71_2_groupi_n_101 = ~(csa_tree_add_71_2_groupi_n_79 & ~csa_tree_add_71_2_groupi_n_97);
 assign csa_tree_add_71_2_groupi_n_100 = ~(csa_tree_add_71_2_groupi_n_75 & (csa_tree_add_71_2_groupi_n_77
    & csa_tree_add_71_2_groupi_n_97));
 assign csa_tree_add_71_2_groupi_n_99 = ~csa_tree_add_71_2_groupi_n_98;
 assign csa_tree_add_71_2_groupi_n_98 = ~(csa_tree_add_71_2_groupi_n_63 & (csa_tree_add_71_2_groupi_n_92
    | csa_tree_add_71_2_groupi_n_68));
 assign csa_tree_add_71_2_groupi_n_97 = ~csa_tree_add_71_2_groupi_n_96;
 assign csa_tree_add_71_2_groupi_n_96 = ~(csa_tree_add_71_2_groupi_n_59 & (csa_tree_add_71_2_groupi_n_58
    & csa_tree_add_71_2_groupi_n_66));
 assign csa_tree_add_71_2_groupi_n_95 = ~(csa_tree_add_71_2_groupi_n_90 | (csa_tree_add_71_2_groupi_n_91
    & csa_tree_add_71_2_groupi_n_83));
 assign csa_tree_add_71_2_groupi_n_94 = ~(csa_tree_add_71_2_groupi_n_82 & csa_tree_add_71_2_groupi_n_67);
 assign csa_tree_add_71_2_groupi_n_93 = ~(csa_tree_add_71_2_groupi_n_82 & csa_tree_add_71_2_groupi_n_83);
 assign csa_tree_add_71_2_groupi_n_91 = ~csa_tree_add_71_2_groupi_n_92;
 assign csa_tree_add_71_2_groupi_n_92 = ~(csa_tree_add_71_2_groupi_n_80 | csa_tree_add_71_2_groupi_n_49);
 assign csa_tree_add_71_2_groupi_n_90 = ~(csa_tree_add_71_2_groupi_n_65 & (csa_tree_add_71_2_groupi_n_60
    | csa_tree_add_71_2_groupi_n_63));
 assign csa_tree_add_71_2_groupi_n_89 = ~(csa_tree_add_71_2_groupi_n_78 & (csa_tree_add_71_2_groupi_n_69
    | csa_tree_add_71_2_groupi_n_64));
 assign csa_tree_add_71_2_groupi_n_88 = ~(csa_tree_add_71_2_groupi_n_67 & csa_tree_add_71_2_groupi_n_63);
 assign csa_tree_add_71_2_groupi_n_87 = ~(csa_tree_add_71_2_groupi_n_70 & csa_tree_add_71_2_groupi_n_78);
 assign csa_tree_add_71_2_groupi_n_81 = ~csa_tree_add_71_2_groupi_n_82;
 assign csa_tree_add_71_2_groupi_n_80 = ~(csa_tree_add_71_2_groupi_n_61 | csa_tree_add_71_2_groupi_n_62);
 assign csa_tree_add_71_2_groupi_n_79 = ~(csa_tree_add_71_2_groupi_n_75 & csa_tree_add_71_2_groupi_n_77);
 assign csa_tree_add_71_2_groupi_n_83 = ~(csa_tree_add_71_2_groupi_n_68 | csa_tree_add_71_2_groupi_n_60);
 assign csa_tree_add_71_2_groupi_n_82 = ~(csa_tree_add_71_2_groupi_n_73 | csa_tree_add_71_2_groupi_n_61);
 assign csa_tree_add_71_2_groupi_n_77 = ~csa_tree_add_71_2_groupi_n_76;
 assign csa_tree_add_71_2_groupi_n_75 = ~csa_tree_add_71_2_groupi_n_74;
 assign csa_tree_add_71_2_groupi_n_72 = ~csa_tree_add_71_2_groupi_n_71;
 assign csa_tree_add_71_2_groupi_n_70 = ~csa_tree_add_71_2_groupi_n_69;
 assign csa_tree_add_71_2_groupi_n_67 = ~csa_tree_add_71_2_groupi_n_68;
 assign csa_tree_add_71_2_groupi_n_66 = ~({in1[0]} & {in3[0]});
 assign csa_tree_add_71_2_groupi_n_78 = ~(csa_tree_add_71_2_groupi_n_3 & csa_tree_add_71_2_groupi_n_9);
 assign csa_tree_add_71_2_groupi_n_76 = (csa_tree_add_71_2_groupi_n_1 & {in3[1]});
 assign csa_tree_add_71_2_groupi_n_74 = ~(csa_tree_add_71_2_groupi_n_1 | {in3[1]});
 assign csa_tree_add_71_2_groupi_n_73 = ~(csa_tree_add_71_2_groupi_n_56 | csa_tree_add_71_2_groupi_n_10);
 assign csa_tree_add_71_2_groupi_n_71 = ~(csa_tree_add_71_2_groupi_n_2 | csa_tree_add_71_2_groupi_n_8);
 assign csa_tree_add_71_2_groupi_n_69 = ~(csa_tree_add_71_2_groupi_n_3 | csa_tree_add_71_2_groupi_n_9);
 assign csa_tree_add_71_2_groupi_n_68 = ~(csa_tree_add_71_2_groupi_n_6 | csa_tree_add_71_2_groupi_n_12);
 assign csa_tree_add_71_2_groupi_n_59 = ~({in1[0]} & {in2[0]});
 assign csa_tree_add_71_2_groupi_n_58 = ~({in3[0]} & {in2[0]});
 assign csa_tree_add_71_2_groupi_n_12 = (({in3[5]} & {in1[5]}) | (({in1[5]} & {in2[5]}) | ({in2[5]} &
    {in3[5]})));
 assign csa_tree_add_71_2_groupi_n_5 = ({in1[5]} ^ ({in2[5]} ^ {in3[5]}));
 assign csa_tree_add_71_2_groupi_n_10 = (({in3[3]} & {in1[3]}) | (({in1[3]} & {in2[3]}) | ({in2[3]} &
    {in3[3]})));
 assign csa_tree_add_71_2_groupi_n_3 = ({in1[3]} ^ ({in2[3]} ^ {in3[3]}));
 assign csa_tree_add_71_2_groupi_n_9 = (({in3[2]} & {in1[2]}) | (({in1[2]} & {in2[2]}) | ({in2[2]} &
    {in3[2]})));
 assign csa_tree_add_71_2_groupi_n_2 = ({in1[2]} ^ ({in2[2]} ^ {in3[2]}));
 assign csa_tree_add_71_2_groupi_n_11 = (({in1[4]} & {in2[4]}) | (({in2[4]} & {in3[4]}) | ({in3[4]} &
    {in1[4]})));
 assign csa_tree_add_71_2_groupi_n_4 = ({in2[4]} ^ ({in3[4]} ^ {in1[4]}));
 assign csa_tree_add_71_2_groupi_n_13 = (({in1[6]} & {in2[6]}) | (({in2[6]} & {in3[6]}) | ({in3[6]} &
    {in1[6]})));
 assign csa_tree_add_71_2_groupi_n_6 = ({in2[6]} ^ ({in3[6]} ^ {in1[6]}));
 assign csa_tree_add_71_2_groupi_n_14 = (({in1[7]} & {in2[7]}) | (({in2[7]} & {in3[7]}) | ({in3[7]} &
    {in1[7]})));
 assign csa_tree_add_71_2_groupi_n_7 = ({in2[7]} ^ ({in3[7]} ^ {in1[7]}));
 assign csa_tree_add_71_2_groupi_n_8 = ({in2[1]} & {in1[1]});
 assign csa_tree_add_71_2_groupi_n_1 = ({in2[1]} ^ {in1[1]});
 assign csa_tree_add_71_2_groupi_n_65 = ~(csa_tree_add_71_2_groupi_n_7 & csa_tree_add_71_2_groupi_n_13);
 assign csa_tree_add_71_2_groupi_n_64 = ~(csa_tree_add_71_2_groupi_n_2 & csa_tree_add_71_2_groupi_n_8);
 assign csa_tree_add_71_2_groupi_n_63 = ~(csa_tree_add_71_2_groupi_n_6 & csa_tree_add_71_2_groupi_n_12);
 assign csa_tree_add_71_2_groupi_n_62 = ~(csa_tree_add_71_2_groupi_n_4 & csa_tree_add_71_2_groupi_n_10);
 assign csa_tree_add_71_2_groupi_n_61 = ~(csa_tree_add_71_2_groupi_n_5 | csa_tree_add_71_2_groupi_n_11);
 assign csa_tree_add_71_2_groupi_n_60 = ~(csa_tree_add_71_2_groupi_n_7 | csa_tree_add_71_2_groupi_n_13);
 assign csa_tree_add_71_2_groupi_n_54 = (csa_tree_add_71_2_groupi_n_61 | csa_tree_add_71_2_groupi_n_49);
 assign csa_tree_add_71_2_groupi_n_53 = ~(csa_tree_add_71_2_groupi_n_60 | ~csa_tree_add_71_2_groupi_n_65);
 assign csa_tree_add_71_2_groupi_n_52 = ~(csa_tree_add_71_2_groupi_n_73 | ~csa_tree_add_71_2_groupi_n_62);
 assign csa_tree_add_71_2_groupi_n_49 = (csa_tree_add_71_2_groupi_n_5 & csa_tree_add_71_2_groupi_n_11);
 assign n_1361 = ((csa_tree_add_86_2_n_982 & csa_tree_add_86_2_n_973) | ((csa_tree_add_86_2_n_973 & csa_tree_add_86_2_n_961)
    | (csa_tree_add_86_2_n_961 & csa_tree_add_86_2_n_982)));
 assign n_1393 = (csa_tree_add_86_2_n_973 ^ (csa_tree_add_86_2_n_961 ^ csa_tree_add_86_2_n_982));
 assign n_1362 = ((csa_tree_add_86_2_n_983 & csa_tree_add_86_2_n_953) | ((csa_tree_add_86_2_n_953 & csa_tree_add_86_2_n_968)
    | (csa_tree_add_86_2_n_968 & csa_tree_add_86_2_n_983)));
 assign n_1394 = (csa_tree_add_86_2_n_953 ^ (csa_tree_add_86_2_n_968 ^ csa_tree_add_86_2_n_983));
 assign n_1360 = ((csa_tree_add_86_2_n_972 & csa_tree_add_86_2_n_945) | ((csa_tree_add_86_2_n_945 & csa_tree_add_86_2_n_960)
    | (csa_tree_add_86_2_n_960 & csa_tree_add_86_2_n_972)));
 assign n_1392 = (csa_tree_add_86_2_n_945 ^ (csa_tree_add_86_2_n_960 ^ csa_tree_add_86_2_n_972));
 assign n_1363 = ((csa_tree_add_86_2_n_974 & csa_tree_add_86_2_n_969) | ((csa_tree_add_86_2_n_969 & csa_tree_add_86_2_n_971)
    | (csa_tree_add_86_2_n_971 & csa_tree_add_86_2_n_974)));
 assign n_1395 = (csa_tree_add_86_2_n_969 ^ (csa_tree_add_86_2_n_971 ^ csa_tree_add_86_2_n_974));
 assign csa_tree_add_86_2_n_982 = ((csa_tree_add_86_2_n_970 & csa_tree_add_86_2_n_899) | ((csa_tree_add_86_2_n_899
    & csa_tree_add_86_2_n_938) | (csa_tree_add_86_2_n_938 & csa_tree_add_86_2_n_970)));
 assign csa_tree_add_86_2_n_983 = (csa_tree_add_86_2_n_899 ^ (csa_tree_add_86_2_n_938 ^ csa_tree_add_86_2_n_970));
 assign n_1364 = ((csa_tree_add_86_2_n_975 & csa_tree_add_86_2_n_947) | ((csa_tree_add_86_2_n_947 & csa_tree_add_86_2_n_954)
    | (csa_tree_add_86_2_n_954 & csa_tree_add_86_2_n_975)));
 assign n_1396 = (csa_tree_add_86_2_n_947 ^ (csa_tree_add_86_2_n_954 ^ csa_tree_add_86_2_n_975));
 assign n_1365 = ((csa_tree_add_86_2_n_964 & csa_tree_add_86_2_n_955) | ((csa_tree_add_86_2_n_955 & csa_tree_add_86_2_n_957)
    | (csa_tree_add_86_2_n_957 & csa_tree_add_86_2_n_964)));
 assign n_1397 = (csa_tree_add_86_2_n_955 ^ (csa_tree_add_86_2_n_957 ^ csa_tree_add_86_2_n_964));
 assign csa_tree_add_86_2_n_974 = ((csa_tree_add_86_2_n_956 & csa_tree_add_86_2_n_941) | ((csa_tree_add_86_2_n_941
    & csa_tree_add_86_2_n_609) | (csa_tree_add_86_2_n_609 & csa_tree_add_86_2_n_956)));
 assign csa_tree_add_86_2_n_975 = (csa_tree_add_86_2_n_941 ^ (csa_tree_add_86_2_n_609 ^ csa_tree_add_86_2_n_956));
 assign csa_tree_add_86_2_n_972 = ((csa_tree_add_86_2_n_952 & csa_tree_add_86_2_n_915) | ((csa_tree_add_86_2_n_915
    & csa_tree_add_86_2_n_611) | (csa_tree_add_86_2_n_611 & csa_tree_add_86_2_n_952)));
 assign csa_tree_add_86_2_n_973 = (csa_tree_add_86_2_n_915 ^ (csa_tree_add_86_2_n_611 ^ csa_tree_add_86_2_n_952));
 assign csa_tree_add_86_2_n_970 = ((csa_tree_add_86_2_n_940 & csa_tree_add_86_2_n_608) | ((csa_tree_add_86_2_n_608
    & csa_tree_add_86_2_n_873) | (csa_tree_add_86_2_n_873 & csa_tree_add_86_2_n_940)));
 assign csa_tree_add_86_2_n_971 = (csa_tree_add_86_2_n_608 ^ (csa_tree_add_86_2_n_873 ^ csa_tree_add_86_2_n_940));
 assign csa_tree_add_86_2_n_968 = ((csa_tree_add_86_2_n_939 & csa_tree_add_86_2_n_919) | ((csa_tree_add_86_2_n_919
    & csa_tree_add_86_2_n_946) | (csa_tree_add_86_2_n_946 & csa_tree_add_86_2_n_939)));
 assign csa_tree_add_86_2_n_969 = (csa_tree_add_86_2_n_919 ^ (csa_tree_add_86_2_n_946 ^ csa_tree_add_86_2_n_939));
 assign n_1359 = ((csa_tree_add_86_2_n_944 & csa_tree_add_86_2_n_755) | ((csa_tree_add_86_2_n_755 & csa_tree_add_86_2_n_685)
    | (csa_tree_add_86_2_n_685 & csa_tree_add_86_2_n_944)));
 assign n_1391 = (csa_tree_add_86_2_n_755 ^ (csa_tree_add_86_2_n_685 ^ csa_tree_add_86_2_n_944));
 assign csa_tree_add_86_2_n_960 = ((csa_tree_add_86_2_n_932 & csa_tree_add_86_2_n_898) | ((csa_tree_add_86_2_n_898
    & csa_tree_add_86_2_n_463) | (csa_tree_add_86_2_n_463 & csa_tree_add_86_2_n_932)));
 assign csa_tree_add_86_2_n_961 = (csa_tree_add_86_2_n_898 ^ (csa_tree_add_86_2_n_463 ^ csa_tree_add_86_2_n_932));
 assign csa_tree_add_86_2_n_952 = ((csa_tree_add_86_2_n_918 & csa_tree_add_86_2_n_933) | ((csa_tree_add_86_2_n_933
    & csa_tree_add_86_2_n_877) | (csa_tree_add_86_2_n_877 & csa_tree_add_86_2_n_918)));
 assign csa_tree_add_86_2_n_953 = (csa_tree_add_86_2_n_933 ^ (csa_tree_add_86_2_n_877 ^ csa_tree_add_86_2_n_918));
 assign csa_tree_add_86_2_n_946 = ((csa_tree_add_86_2_n_907 & csa_tree_add_86_2_n_912) | ((csa_tree_add_86_2_n_912
    & csa_tree_add_86_2_n_668) | (csa_tree_add_86_2_n_668 & csa_tree_add_86_2_n_907)));
 assign csa_tree_add_86_2_n_947 = (csa_tree_add_86_2_n_912 ^ (csa_tree_add_86_2_n_668 ^ csa_tree_add_86_2_n_907));
 assign csa_tree_add_86_2_n_944 = ((csa_tree_add_86_2_n_914 & csa_tree_add_86_2_n_551) | ((csa_tree_add_86_2_n_551
    & csa_tree_add_86_2_n_703) | (csa_tree_add_86_2_n_703 & csa_tree_add_86_2_n_914)));
 assign csa_tree_add_86_2_n_945 = (csa_tree_add_86_2_n_551 ^ (csa_tree_add_86_2_n_703 ^ csa_tree_add_86_2_n_914));
 assign csa_tree_add_86_2_n_938 = ((csa_tree_add_86_2_n_906 & csa_tree_add_86_2_n_115) | ((csa_tree_add_86_2_n_115
    & csa_tree_add_86_2_n_897) | (csa_tree_add_86_2_n_897 & csa_tree_add_86_2_n_906)));
 assign csa_tree_add_86_2_n_939 = (csa_tree_add_86_2_n_115 ^ (csa_tree_add_86_2_n_897 ^ csa_tree_add_86_2_n_906));
 assign csa_tree_add_86_2_n_932 = ((csa_tree_add_86_2_n_896 & csa_tree_add_86_2_n_103) | ((csa_tree_add_86_2_n_103
    & csa_tree_add_86_2_n_441) | (csa_tree_add_86_2_n_441 & csa_tree_add_86_2_n_896)));
 assign csa_tree_add_86_2_n_933 = (csa_tree_add_86_2_n_103 ^ (csa_tree_add_86_2_n_441 ^ csa_tree_add_86_2_n_896));
 assign csa_tree_add_86_2_n_920 = ((csa_tree_add_86_2_n_892 & csa_tree_add_86_2_n_139) | ((csa_tree_add_86_2_n_139
    & csa_tree_add_86_2_n_875) | (csa_tree_add_86_2_n_875 & csa_tree_add_86_2_n_892)));
 assign csa_tree_add_86_2_n_921 = (csa_tree_add_86_2_n_139 ^ (csa_tree_add_86_2_n_875 ^ csa_tree_add_86_2_n_892));
 assign csa_tree_add_86_2_n_914 = ((csa_tree_add_86_2_n_876 & csa_tree_add_86_2_n_138) | ((csa_tree_add_86_2_n_138
    & csa_tree_add_86_2_n_79) | (csa_tree_add_86_2_n_79 & csa_tree_add_86_2_n_876)));
 assign csa_tree_add_86_2_n_915 = (csa_tree_add_86_2_n_138 ^ (csa_tree_add_86_2_n_79 ^ csa_tree_add_86_2_n_876));
 assign n_1370 = ((csa_tree_add_86_2_n_885 & csa_tree_add_86_2_n_837) | ((csa_tree_add_86_2_n_837 & csa_tree_add_86_2_n_834)
    | (csa_tree_add_86_2_n_834 & csa_tree_add_86_2_n_885)));
 assign n_1401 = (csa_tree_add_86_2_n_837 ^ (csa_tree_add_86_2_n_834 ^ csa_tree_add_86_2_n_885));
 assign csa_tree_add_86_2_n_902 = ((csa_tree_add_86_2_n_826 & csa_tree_add_86_2_n_845) | ((csa_tree_add_86_2_n_845
    & csa_tree_add_86_2_n_860) | (csa_tree_add_86_2_n_860 & csa_tree_add_86_2_n_826)));
 assign csa_tree_add_86_2_n_903 = (csa_tree_add_86_2_n_845 ^ (csa_tree_add_86_2_n_860 ^ csa_tree_add_86_2_n_826));
 assign csa_tree_add_86_2_n_898 = ((csa_tree_add_86_2_n_872 & csa_tree_add_86_2_n_160) | ((csa_tree_add_86_2_n_160
    & csa_tree_add_86_2_n_163) | (csa_tree_add_86_2_n_163 & csa_tree_add_86_2_n_872)));
 assign csa_tree_add_86_2_n_899 = (csa_tree_add_86_2_n_160 ^ (csa_tree_add_86_2_n_163 ^ csa_tree_add_86_2_n_872));
 assign csa_tree_add_86_2_n_894 = ((csa_tree_add_86_2_n_851 & csa_tree_add_86_2_n_836) | ((csa_tree_add_86_2_n_836
    & csa_tree_add_86_2_n_839) | (csa_tree_add_86_2_n_839 & csa_tree_add_86_2_n_851)));
 assign csa_tree_add_86_2_n_895 = (csa_tree_add_86_2_n_836 ^ (csa_tree_add_86_2_n_839 ^ csa_tree_add_86_2_n_851));
 assign csa_tree_add_86_2_n_892 = ((csa_tree_add_86_2_n_861 & csa_tree_add_86_2_n_74) | ((csa_tree_add_86_2_n_74
    & csa_tree_add_86_2_n_842) | (csa_tree_add_86_2_n_842 & csa_tree_add_86_2_n_861)));
 assign csa_tree_add_86_2_n_893 = (csa_tree_add_86_2_n_74 ^ (csa_tree_add_86_2_n_842 ^ csa_tree_add_86_2_n_861));
 assign csa_tree_add_86_2_n_890 = ((csa_tree_add_86_2_n_854 & csa_tree_add_86_2_n_141) | ((csa_tree_add_86_2_n_141
    & csa_tree_add_86_2_n_840) | (csa_tree_add_86_2_n_840 & csa_tree_add_86_2_n_854)));
 assign csa_tree_add_86_2_n_891 = (csa_tree_add_86_2_n_141 ^ (csa_tree_add_86_2_n_840 ^ csa_tree_add_86_2_n_854));
 assign csa_tree_add_86_2_n_888 = ((csa_tree_add_86_2_n_852 & csa_tree_add_86_2_n_52) | ((csa_tree_add_86_2_n_52
    & csa_tree_add_86_2_n_843) | (csa_tree_add_86_2_n_843 & csa_tree_add_86_2_n_852)));
 assign csa_tree_add_86_2_n_889 = (csa_tree_add_86_2_n_52 ^ (csa_tree_add_86_2_n_843 ^ csa_tree_add_86_2_n_852));
 assign csa_tree_add_86_2_n_886 = ((csa_tree_add_86_2_n_853 & csa_tree_add_86_2_n_98) | ((csa_tree_add_86_2_n_98
    & csa_tree_add_86_2_n_850) | (csa_tree_add_86_2_n_850 & csa_tree_add_86_2_n_853)));
 assign csa_tree_add_86_2_n_887 = (csa_tree_add_86_2_n_98 ^ (csa_tree_add_86_2_n_850 ^ csa_tree_add_86_2_n_853));
 assign csa_tree_add_86_2_n_884 = ((csa_tree_add_86_2_n_849 & csa_tree_add_86_2_n_785) | ((csa_tree_add_86_2_n_785
    & csa_tree_add_86_2_n_824) | (csa_tree_add_86_2_n_824 & csa_tree_add_86_2_n_849)));
 assign csa_tree_add_86_2_n_885 = (csa_tree_add_86_2_n_785 ^ (csa_tree_add_86_2_n_824 ^ csa_tree_add_86_2_n_849));
 assign csa_tree_add_86_2_n_882 = ((csa_tree_add_86_2_n_841 & csa_tree_add_86_2_n_83) | ((csa_tree_add_86_2_n_83
    & csa_tree_add_86_2_n_41) | (csa_tree_add_86_2_n_41 & csa_tree_add_86_2_n_841)));
 assign csa_tree_add_86_2_n_883 = (csa_tree_add_86_2_n_83 ^ (csa_tree_add_86_2_n_41 ^ csa_tree_add_86_2_n_841));
 assign csa_tree_add_86_2_n_874 = ((csa_tree_add_86_2_n_831 & csa_tree_add_86_2_n_188) | ((csa_tree_add_86_2_n_188
    & csa_tree_add_86_2_n_814) | (csa_tree_add_86_2_n_814 & csa_tree_add_86_2_n_831)));
 assign csa_tree_add_86_2_n_875 = (csa_tree_add_86_2_n_188 ^ (csa_tree_add_86_2_n_814 ^ csa_tree_add_86_2_n_831));
 assign csa_tree_add_86_2_n_870 = ((csa_tree_add_86_2_n_827 & csa_tree_add_86_2_n_186) | ((csa_tree_add_86_2_n_186
    & csa_tree_add_86_2_n_151) | (csa_tree_add_86_2_n_151 & csa_tree_add_86_2_n_827)));
 assign csa_tree_add_86_2_n_871 = (csa_tree_add_86_2_n_186 ^ (csa_tree_add_86_2_n_151 ^ csa_tree_add_86_2_n_827));
 assign csa_tree_add_86_2_n_868 = ((csa_tree_add_86_2_n_848 & csa_tree_add_86_2_n_66) | ((csa_tree_add_86_2_n_66
    & csa_tree_add_86_2_n_803) | (csa_tree_add_86_2_n_803 & csa_tree_add_86_2_n_848)));
 assign csa_tree_add_86_2_n_869 = (csa_tree_add_86_2_n_66 ^ (csa_tree_add_86_2_n_803 ^ csa_tree_add_86_2_n_848));
 assign n_1371 = ((csa_tree_add_86_2_n_835 & csa_tree_add_86_2_n_764) | ((csa_tree_add_86_2_n_764 & csa_tree_add_86_2_n_825)
    | (csa_tree_add_86_2_n_825 & csa_tree_add_86_2_n_835)));
 assign n_1402 = (csa_tree_add_86_2_n_764 ^ (csa_tree_add_86_2_n_825 ^ csa_tree_add_86_2_n_835));
 assign csa_tree_add_86_2_n_862 = ((csa_tree_add_86_2_n_838 & csa_tree_add_86_2_n_166) | ((csa_tree_add_86_2_n_166
    & csa_tree_add_86_2_n_821) | (csa_tree_add_86_2_n_821 & csa_tree_add_86_2_n_838)));
 assign csa_tree_add_86_2_n_863 = (csa_tree_add_86_2_n_166 ^ (csa_tree_add_86_2_n_821 ^ csa_tree_add_86_2_n_838));
 assign csa_tree_add_86_2_n_860 = ((csa_tree_add_86_2_n_790 & csa_tree_add_86_2_n_774) | ((csa_tree_add_86_2_n_774
    & csa_tree_add_86_2_n_817) | (csa_tree_add_86_2_n_817 & csa_tree_add_86_2_n_790)));
 assign csa_tree_add_86_2_n_861 = (csa_tree_add_86_2_n_774 ^ (csa_tree_add_86_2_n_817 ^ csa_tree_add_86_2_n_790));
 assign csa_tree_add_86_2_n_858 = ((csa_tree_add_86_2_n_802 & csa_tree_add_86_2_n_164) | ((csa_tree_add_86_2_n_164
    & csa_tree_add_86_2_n_804) | (csa_tree_add_86_2_n_804 & csa_tree_add_86_2_n_802)));
 assign csa_tree_add_86_2_n_859 = (csa_tree_add_86_2_n_164 ^ (csa_tree_add_86_2_n_804 ^ csa_tree_add_86_2_n_802));
 assign csa_tree_add_86_2_n_854 = ((csa_tree_add_86_2_n_791 & csa_tree_add_86_2_n_173) | ((csa_tree_add_86_2_n_173
    & csa_tree_add_86_2_n_820) | (csa_tree_add_86_2_n_820 & csa_tree_add_86_2_n_791)));
 assign csa_tree_add_86_2_n_855 = (csa_tree_add_86_2_n_173 ^ (csa_tree_add_86_2_n_820 ^ csa_tree_add_86_2_n_791));
 assign csa_tree_add_86_2_n_852 = ((csa_tree_add_86_2_n_807 & csa_tree_add_86_2_n_47) | ((csa_tree_add_86_2_n_47
    & csa_tree_add_86_2_n_789) | (csa_tree_add_86_2_n_789 & csa_tree_add_86_2_n_807)));
 assign csa_tree_add_86_2_n_853 = (csa_tree_add_86_2_n_47 ^ (csa_tree_add_86_2_n_789 ^ csa_tree_add_86_2_n_807));
 assign csa_tree_add_86_2_n_850 = ((csa_tree_add_86_2_n_805 & csa_tree_add_86_2_n_76) | ((csa_tree_add_86_2_n_76
    & csa_tree_add_86_2_n_106) | (csa_tree_add_86_2_n_106 & csa_tree_add_86_2_n_805)));
 assign csa_tree_add_86_2_n_851 = (csa_tree_add_86_2_n_76 ^ (csa_tree_add_86_2_n_106 ^ csa_tree_add_86_2_n_805));
 assign csa_tree_add_86_2_n_848 = ((csa_tree_add_86_2_n_780 & csa_tree_add_86_2_n_86) | ((csa_tree_add_86_2_n_86
    & csa_tree_add_86_2_n_782) | (csa_tree_add_86_2_n_782 & csa_tree_add_86_2_n_780)));
 assign csa_tree_add_86_2_n_849 = (csa_tree_add_86_2_n_86 ^ (csa_tree_add_86_2_n_782 ^ csa_tree_add_86_2_n_780));
 assign n_1372 = ((csa_tree_add_86_2_n_776 & csa_tree_add_86_2_n_742) | ((csa_tree_add_86_2_n_742 & csa_tree_add_86_2_n_779)
    | (csa_tree_add_86_2_n_779 & csa_tree_add_86_2_n_776)));
 assign n_1403 = (csa_tree_add_86_2_n_742 ^ (csa_tree_add_86_2_n_779 ^ csa_tree_add_86_2_n_776));
 assign csa_tree_add_86_2_n_844 = ((csa_tree_add_86_2_n_799 & csa_tree_add_86_2_n_54) | ((csa_tree_add_86_2_n_54
    & csa_tree_add_86_2_n_222) | (csa_tree_add_86_2_n_222 & csa_tree_add_86_2_n_799)));
 assign csa_tree_add_86_2_n_845 = (csa_tree_add_86_2_n_54 ^ (csa_tree_add_86_2_n_222 ^ csa_tree_add_86_2_n_799));
 assign csa_tree_add_86_2_n_842 = ((csa_tree_add_86_2_n_788 & csa_tree_add_86_2_n_162) | ((csa_tree_add_86_2_n_162
    & csa_tree_add_86_2_n_737) | (csa_tree_add_86_2_n_737 & csa_tree_add_86_2_n_788)));
 assign csa_tree_add_86_2_n_843 = (csa_tree_add_86_2_n_162 ^ (csa_tree_add_86_2_n_737 ^ csa_tree_add_86_2_n_788));
 assign csa_tree_add_86_2_n_840 = ((csa_tree_add_86_2_n_806 & csa_tree_add_86_2_n_42) | ((csa_tree_add_86_2_n_42
    & csa_tree_add_86_2_n_775) | (csa_tree_add_86_2_n_775 & csa_tree_add_86_2_n_806)));
 assign csa_tree_add_86_2_n_841 = (csa_tree_add_86_2_n_42 ^ (csa_tree_add_86_2_n_775 ^ csa_tree_add_86_2_n_806));
 assign csa_tree_add_86_2_n_838 = ((csa_tree_add_86_2_n_784 & csa_tree_add_86_2_n_157) | ((csa_tree_add_86_2_n_157
    & csa_tree_add_86_2_n_768) | (csa_tree_add_86_2_n_768 & csa_tree_add_86_2_n_784)));
 assign csa_tree_add_86_2_n_839 = (csa_tree_add_86_2_n_157 ^ (csa_tree_add_86_2_n_768 ^ csa_tree_add_86_2_n_784));
 assign csa_tree_add_86_2_n_836 = ((csa_tree_add_86_2_n_769 & csa_tree_add_86_2_n_67) | ((csa_tree_add_86_2_n_67
    & csa_tree_add_86_2_n_101) | (csa_tree_add_86_2_n_101 & csa_tree_add_86_2_n_769)));
 assign csa_tree_add_86_2_n_837 = (csa_tree_add_86_2_n_67 ^ (csa_tree_add_86_2_n_101 ^ csa_tree_add_86_2_n_769));
 assign csa_tree_add_86_2_n_834 = ((csa_tree_add_86_2_n_781 & csa_tree_add_86_2_n_131) | ((csa_tree_add_86_2_n_131
    & csa_tree_add_86_2_n_778) | (csa_tree_add_86_2_n_778 & csa_tree_add_86_2_n_781)));
 assign csa_tree_add_86_2_n_835 = (csa_tree_add_86_2_n_131 ^ (csa_tree_add_86_2_n_778 ^ csa_tree_add_86_2_n_781));
 assign csa_tree_add_86_2_n_832 = ((csa_tree_add_86_2_n_798 & csa_tree_add_86_2_n_699) | ((csa_tree_add_86_2_n_699
    & csa_tree_add_86_2_n_759) | (csa_tree_add_86_2_n_759 & csa_tree_add_86_2_n_798)));
 assign csa_tree_add_86_2_n_833 = (csa_tree_add_86_2_n_699 ^ (csa_tree_add_86_2_n_759 ^ csa_tree_add_86_2_n_798));
 assign csa_tree_add_86_2_n_830 = ((csa_tree_add_86_2_n_816 & csa_tree_add_86_2_n_238) | ((csa_tree_add_86_2_n_238
    & csa_tree_add_86_2_n_756) | (csa_tree_add_86_2_n_756 & csa_tree_add_86_2_n_816)));
 assign csa_tree_add_86_2_n_831 = (csa_tree_add_86_2_n_238 ^ (csa_tree_add_86_2_n_756 ^ csa_tree_add_86_2_n_816));
 assign csa_tree_add_86_2_n_826 = ((csa_tree_add_86_2_n_815 & csa_tree_add_86_2_n_81) | ((csa_tree_add_86_2_n_81
    & csa_tree_add_86_2_n_111) | (csa_tree_add_86_2_n_111 & csa_tree_add_86_2_n_815)));
 assign csa_tree_add_86_2_n_827 = (csa_tree_add_86_2_n_81 ^ (csa_tree_add_86_2_n_111 ^ csa_tree_add_86_2_n_815));
 assign csa_tree_add_86_2_n_824 = ((csa_tree_add_86_2_n_783 & csa_tree_add_86_2_n_61) | ((csa_tree_add_86_2_n_61
    & csa_tree_add_86_2_n_147) | (csa_tree_add_86_2_n_147 & csa_tree_add_86_2_n_783)));
 assign csa_tree_add_86_2_n_825 = (csa_tree_add_86_2_n_61 ^ (csa_tree_add_86_2_n_147 ^ csa_tree_add_86_2_n_783));
 assign n_1358 = ((csa_tree_add_86_2_n_723 & csa_tree_add_86_2_n_754) | ((csa_tree_add_86_2_n_754 & csa_tree_add_86_2_n_684)
    | (csa_tree_add_86_2_n_684 & csa_tree_add_86_2_n_723)));
 assign n_1390 = (csa_tree_add_86_2_n_754 ^ (csa_tree_add_86_2_n_684 ^ csa_tree_add_86_2_n_723));
 assign csa_tree_add_86_2_n_820 = ((csa_tree_add_86_2_n_719 & csa_tree_add_86_2_n_175) | ((csa_tree_add_86_2_n_175
    & csa_tree_add_86_2_n_760) | (csa_tree_add_86_2_n_760 & csa_tree_add_86_2_n_719)));
 assign csa_tree_add_86_2_n_821 = (csa_tree_add_86_2_n_175 ^ (csa_tree_add_86_2_n_760 ^ csa_tree_add_86_2_n_719));
 assign csa_tree_add_86_2_n_818 = ((csa_tree_add_86_2_n_758 & csa_tree_add_86_2_n_698) | ((csa_tree_add_86_2_n_698
    & csa_tree_add_86_2_n_753) | (csa_tree_add_86_2_n_753 & csa_tree_add_86_2_n_758)));
 assign csa_tree_add_86_2_n_819 = (csa_tree_add_86_2_n_698 ^ (csa_tree_add_86_2_n_753 ^ csa_tree_add_86_2_n_758));
 assign csa_tree_add_86_2_n_816 = ((csa_tree_add_86_2_n_736 & csa_tree_add_86_2_n_738) | ((csa_tree_add_86_2_n_738
    & csa_tree_add_86_2_n_747) | (csa_tree_add_86_2_n_747 & csa_tree_add_86_2_n_736)));
 assign csa_tree_add_86_2_n_817 = (csa_tree_add_86_2_n_738 ^ (csa_tree_add_86_2_n_747 ^ csa_tree_add_86_2_n_736));
 assign csa_tree_add_86_2_n_814 = ((csa_tree_add_86_2_n_757 & csa_tree_add_86_2_n_169) | ((csa_tree_add_86_2_n_169
    & csa_tree_add_86_2_n_229) | (csa_tree_add_86_2_n_229 & csa_tree_add_86_2_n_757)));
 assign csa_tree_add_86_2_n_815 = (csa_tree_add_86_2_n_169 ^ (csa_tree_add_86_2_n_229 ^ csa_tree_add_86_2_n_757));
 assign n_1357 = ((csa_tree_add_86_2_n_722 & csa_tree_add_86_2_n_745) | ((csa_tree_add_86_2_n_745 & csa_tree_add_86_2_n_689)
    | (csa_tree_add_86_2_n_689 & csa_tree_add_86_2_n_722)));
 assign n_1389 = (csa_tree_add_86_2_n_745 ^ (csa_tree_add_86_2_n_689 ^ csa_tree_add_86_2_n_722));
 assign n_1353 = ((csa_tree_add_86_2_n_732 & csa_tree_add_86_2_n_735) | ((csa_tree_add_86_2_n_735 & csa_tree_add_86_2_n_687)
    | (csa_tree_add_86_2_n_687 & csa_tree_add_86_2_n_732)));
 assign n_1385 = (csa_tree_add_86_2_n_735 ^ (csa_tree_add_86_2_n_687 ^ csa_tree_add_86_2_n_732));
 assign csa_tree_add_86_2_n_806 = ((csa_tree_add_86_2_n_751 & csa_tree_add_86_2_n_122) | ((csa_tree_add_86_2_n_122
    & csa_tree_add_86_2_n_694) | (csa_tree_add_86_2_n_694 & csa_tree_add_86_2_n_751)));
 assign csa_tree_add_86_2_n_807 = (csa_tree_add_86_2_n_122 ^ (csa_tree_add_86_2_n_694 ^ csa_tree_add_86_2_n_751));
 assign csa_tree_add_86_2_n_804 = ((csa_tree_add_86_2_n_748 & csa_tree_add_86_2_n_714) | ((csa_tree_add_86_2_n_714
    & csa_tree_add_86_2_n_731) | (csa_tree_add_86_2_n_731 & csa_tree_add_86_2_n_748)));
 assign csa_tree_add_86_2_n_805 = (csa_tree_add_86_2_n_714 ^ (csa_tree_add_86_2_n_731 ^ csa_tree_add_86_2_n_748));
 assign csa_tree_add_86_2_n_802 = ((csa_tree_add_86_2_n_761 & csa_tree_add_86_2_n_68) | ((csa_tree_add_86_2_n_68
    & csa_tree_add_86_2_n_695) | (csa_tree_add_86_2_n_695 & csa_tree_add_86_2_n_761)));
 assign csa_tree_add_86_2_n_803 = (csa_tree_add_86_2_n_68 ^ (csa_tree_add_86_2_n_695 ^ csa_tree_add_86_2_n_761));
 assign n_1356 = ((csa_tree_add_86_2_n_744 & csa_tree_add_86_2_n_727) | ((csa_tree_add_86_2_n_727 & csa_tree_add_86_2_n_688)
    | (csa_tree_add_86_2_n_688 & csa_tree_add_86_2_n_744)));
 assign n_1388 = (csa_tree_add_86_2_n_727 ^ (csa_tree_add_86_2_n_688 ^ csa_tree_add_86_2_n_744));
 assign csa_tree_add_86_2_n_798 = ((csa_tree_add_86_2_n_746 & csa_tree_add_86_2_n_725) | ((csa_tree_add_86_2_n_725
    & csa_tree_add_86_2_n_647) | (csa_tree_add_86_2_n_647 & csa_tree_add_86_2_n_746)));
 assign csa_tree_add_86_2_n_799 = (csa_tree_add_86_2_n_725 ^ (csa_tree_add_86_2_n_647 ^ csa_tree_add_86_2_n_746));
 assign csa_tree_add_86_2_n_790 = ((csa_tree_add_86_2_n_739 & csa_tree_add_86_2_n_127) | ((csa_tree_add_86_2_n_127
    & csa_tree_add_86_2_n_718) | (csa_tree_add_86_2_n_718 & csa_tree_add_86_2_n_739)));
 assign csa_tree_add_86_2_n_791 = (csa_tree_add_86_2_n_127 ^ (csa_tree_add_86_2_n_718 ^ csa_tree_add_86_2_n_739));
 assign csa_tree_add_86_2_n_788 = ((csa_tree_add_86_2_n_730 & csa_tree_add_86_2_n_161) | ((csa_tree_add_86_2_n_161
    & csa_tree_add_86_2_n_701) | (csa_tree_add_86_2_n_701 & csa_tree_add_86_2_n_730)));
 assign csa_tree_add_86_2_n_789 = (csa_tree_add_86_2_n_161 ^ (csa_tree_add_86_2_n_701 ^ csa_tree_add_86_2_n_730));
 assign n_1355 = ((csa_tree_add_86_2_n_726 & csa_tree_add_86_2_n_717) | ((csa_tree_add_86_2_n_717 & csa_tree_add_86_2_n_679)
    | (csa_tree_add_86_2_n_679 & csa_tree_add_86_2_n_726)));
 assign n_1387 = (csa_tree_add_86_2_n_717 ^ (csa_tree_add_86_2_n_679 ^ csa_tree_add_86_2_n_726));
 assign csa_tree_add_86_2_n_784 = ((csa_tree_add_86_2_n_749 & csa_tree_add_86_2_n_57) | ((csa_tree_add_86_2_n_57
    & csa_tree_add_86_2_n_712) | (csa_tree_add_86_2_n_712 & csa_tree_add_86_2_n_749)));
 assign csa_tree_add_86_2_n_785 = (csa_tree_add_86_2_n_57 ^ (csa_tree_add_86_2_n_712 ^ csa_tree_add_86_2_n_749));
 assign csa_tree_add_86_2_n_782 = ((csa_tree_add_86_2_n_675 & csa_tree_add_86_2_n_82) | ((csa_tree_add_86_2_n_82
    & csa_tree_add_86_2_n_690) | (csa_tree_add_86_2_n_690 & csa_tree_add_86_2_n_675)));
 assign csa_tree_add_86_2_n_783 = (csa_tree_add_86_2_n_82 ^ (csa_tree_add_86_2_n_690 ^ csa_tree_add_86_2_n_675));
 assign csa_tree_add_86_2_n_780 = ((csa_tree_add_86_2_n_713 & csa_tree_add_86_2_n_59) | ((csa_tree_add_86_2_n_59
    & csa_tree_add_86_2_n_710) | (csa_tree_add_86_2_n_710 & csa_tree_add_86_2_n_713)));
 assign csa_tree_add_86_2_n_781 = (csa_tree_add_86_2_n_59 ^ (csa_tree_add_86_2_n_710 ^ csa_tree_add_86_2_n_713));
 assign csa_tree_add_86_2_n_778 = ((csa_tree_add_86_2_n_708 & csa_tree_add_86_2_n_75) | ((csa_tree_add_86_2_n_75
    & csa_tree_add_86_2_n_691) | (csa_tree_add_86_2_n_691 & csa_tree_add_86_2_n_708)));
 assign csa_tree_add_86_2_n_779 = (csa_tree_add_86_2_n_75 ^ (csa_tree_add_86_2_n_691 ^ csa_tree_add_86_2_n_708));
 assign csa_tree_add_86_2_n_776 = ((csa_tree_add_86_2_n_706 & csa_tree_add_86_2_n_179) | ((csa_tree_add_86_2_n_179
    & csa_tree_add_86_2_n_709) | (csa_tree_add_86_2_n_709 & csa_tree_add_86_2_n_706)));
 assign n_1404 = (csa_tree_add_86_2_n_179 ^ (csa_tree_add_86_2_n_709 ^ csa_tree_add_86_2_n_706));
 assign csa_tree_add_86_2_n_774 = ((csa_tree_add_86_2_n_750 & csa_tree_add_86_2_n_231) | ((csa_tree_add_86_2_n_231
    & csa_tree_add_86_2_n_700) | (csa_tree_add_86_2_n_700 & csa_tree_add_86_2_n_750)));
 assign csa_tree_add_86_2_n_775 = (csa_tree_add_86_2_n_231 ^ (csa_tree_add_86_2_n_700 ^ csa_tree_add_86_2_n_750));
 assign csa_tree_add_86_2_n_772 = ((csa_tree_add_86_2_n_752 & csa_tree_add_86_2_n_652) | ((csa_tree_add_86_2_n_652
    & csa_tree_add_86_2_n_557) | (csa_tree_add_86_2_n_557 & csa_tree_add_86_2_n_752)));
 assign csa_tree_add_86_2_n_773 = (csa_tree_add_86_2_n_652 ^ (csa_tree_add_86_2_n_557 ^ csa_tree_add_86_2_n_752));
 assign csa_tree_add_86_2_n_768 = ((csa_tree_add_86_2_n_715 & csa_tree_add_86_2_n_44) | ((csa_tree_add_86_2_n_44
    & csa_tree_add_86_2_n_697) | (csa_tree_add_86_2_n_697 & csa_tree_add_86_2_n_715)));
 assign csa_tree_add_86_2_n_769 = (csa_tree_add_86_2_n_44 ^ (csa_tree_add_86_2_n_697 ^ csa_tree_add_86_2_n_715));
 assign n_1354 = ((csa_tree_add_86_2_n_716 & csa_tree_add_86_2_n_733) | ((csa_tree_add_86_2_n_733 & csa_tree_add_86_2_n_681)
    | (csa_tree_add_86_2_n_681 & csa_tree_add_86_2_n_716)));
 assign n_1386 = (csa_tree_add_86_2_n_733 ^ (csa_tree_add_86_2_n_681 ^ csa_tree_add_86_2_n_716));
 assign csa_tree_add_86_2_n_764 = ((csa_tree_add_86_2_n_711 & csa_tree_add_86_2_n_172) | ((csa_tree_add_86_2_n_172
    & csa_tree_add_86_2_n_133) | (csa_tree_add_86_2_n_133 & csa_tree_add_86_2_n_711)));
 assign n_1373 = (csa_tree_add_86_2_n_172 ^ (csa_tree_add_86_2_n_133 ^ csa_tree_add_86_2_n_711));
 assign csa_tree_add_86_2_n_762 = ((csa_tree_add_86_2_n_704 & csa_tree_add_86_2_n_555) | ((csa_tree_add_86_2_n_555
    & csa_tree_add_86_2_n_683) | (csa_tree_add_86_2_n_683 & csa_tree_add_86_2_n_704)));
 assign n_1379 = (csa_tree_add_86_2_n_555 ^ (csa_tree_add_86_2_n_683 ^ csa_tree_add_86_2_n_704));
 assign csa_tree_add_86_2_n_760 = ((csa_tree_add_86_2_n_651 & csa_tree_add_86_2_n_140) | ((csa_tree_add_86_2_n_140
    & csa_tree_add_86_2_n_696) | (csa_tree_add_86_2_n_696 & csa_tree_add_86_2_n_651)));
 assign csa_tree_add_86_2_n_761 = (csa_tree_add_86_2_n_140 ^ (csa_tree_add_86_2_n_696 ^ csa_tree_add_86_2_n_651));
 assign csa_tree_add_86_2_n_758 = ((csa_tree_add_86_2_n_724 & csa_tree_add_86_2_n_646) | ((csa_tree_add_86_2_n_646
    & csa_tree_add_86_2_n_625) | (csa_tree_add_86_2_n_625 & csa_tree_add_86_2_n_724)));
 assign csa_tree_add_86_2_n_759 = (csa_tree_add_86_2_n_646 ^ (csa_tree_add_86_2_n_625 ^ csa_tree_add_86_2_n_724));
 assign csa_tree_add_86_2_n_756 = ((csa_tree_add_86_2_n_663 & csa_tree_add_86_2_n_656) | ((csa_tree_add_86_2_n_656
    & csa_tree_add_86_2_n_659) | (csa_tree_add_86_2_n_659 & csa_tree_add_86_2_n_663)));
 assign csa_tree_add_86_2_n_757 = (csa_tree_add_86_2_n_656 ^ (csa_tree_add_86_2_n_659 ^ csa_tree_add_86_2_n_663));
 assign csa_tree_add_86_2_n_754 = ((csa_tree_add_86_2_n_702 & csa_tree_add_86_2_n_607) | ((csa_tree_add_86_2_n_607
    & csa_tree_add_86_2_n_550) | (csa_tree_add_86_2_n_550 & csa_tree_add_86_2_n_702)));
 assign csa_tree_add_86_2_n_755 = (csa_tree_add_86_2_n_607 ^ (csa_tree_add_86_2_n_550 ^ csa_tree_add_86_2_n_702));
 assign csa_tree_add_86_2_n_752 = ((csa_tree_add_86_2_n_624 & csa_tree_add_86_2_n_467) | ((csa_tree_add_86_2_n_467
    & csa_tree_add_86_2_n_653) | (csa_tree_add_86_2_n_653 & csa_tree_add_86_2_n_624)));
 assign csa_tree_add_86_2_n_753 = (csa_tree_add_86_2_n_467 ^ (csa_tree_add_86_2_n_653 ^ csa_tree_add_86_2_n_624));
 assign csa_tree_add_86_2_n_750 = ((csa_tree_add_86_2_n_631 & csa_tree_add_86_2_n_626) | ((csa_tree_add_86_2_n_626
    & csa_tree_add_86_2_n_655) | (csa_tree_add_86_2_n_655 & csa_tree_add_86_2_n_631)));
 assign csa_tree_add_86_2_n_751 = (csa_tree_add_86_2_n_626 ^ (csa_tree_add_86_2_n_655 ^ csa_tree_add_86_2_n_631));
 assign csa_tree_add_86_2_n_748 = ((csa_tree_add_86_2_n_674 & csa_tree_add_86_2_n_94) | ((csa_tree_add_86_2_n_94
    & csa_tree_add_86_2_n_649) | (csa_tree_add_86_2_n_649 & csa_tree_add_86_2_n_674)));
 assign csa_tree_add_86_2_n_749 = (csa_tree_add_86_2_n_94 ^ (csa_tree_add_86_2_n_649 ^ csa_tree_add_86_2_n_674));
 assign csa_tree_add_86_2_n_746 = ((csa_tree_add_86_2_n_664 & csa_tree_add_86_2_n_638) | ((csa_tree_add_86_2_n_638
    & csa_tree_add_86_2_n_525) | (csa_tree_add_86_2_n_525 & csa_tree_add_86_2_n_664)));
 assign csa_tree_add_86_2_n_747 = (csa_tree_add_86_2_n_638 ^ (csa_tree_add_86_2_n_525 ^ csa_tree_add_86_2_n_664));
 assign csa_tree_add_86_2_n_744 = ((csa_tree_add_86_2_n_670 & csa_tree_add_86_2_n_635) | ((csa_tree_add_86_2_n_635
    & csa_tree_add_86_2_n_561) | (csa_tree_add_86_2_n_561 & csa_tree_add_86_2_n_670)));
 assign csa_tree_add_86_2_n_745 = (csa_tree_add_86_2_n_635 ^ (csa_tree_add_86_2_n_561 ^ csa_tree_add_86_2_n_670));
 assign csa_tree_add_86_2_n_742 = ((csa_tree_add_86_2_n_660 & csa_tree_add_86_2_n_144) | ((csa_tree_add_86_2_n_144
    & csa_tree_add_86_2_n_153) | (csa_tree_add_86_2_n_153 & csa_tree_add_86_2_n_660)));
 assign n_1374 = (csa_tree_add_86_2_n_144 ^ (csa_tree_add_86_2_n_153 ^ csa_tree_add_86_2_n_660));
 assign csa_tree_add_86_2_n_740 = ((csa_tree_add_86_2_n_686 & csa_tree_add_86_2_n_585) | ((csa_tree_add_86_2_n_585
    & csa_tree_add_86_2_n_602) | (csa_tree_add_86_2_n_602 & csa_tree_add_86_2_n_686)));
 assign csa_tree_add_86_2_n_741 = (csa_tree_add_86_2_n_585 ^ (csa_tree_add_86_2_n_602 ^ csa_tree_add_86_2_n_686));
 assign csa_tree_add_86_2_n_738 = ((csa_tree_add_86_2_n_630 & csa_tree_add_86_2_n_654) | ((csa_tree_add_86_2_n_654
    & csa_tree_add_86_2_n_639) | (csa_tree_add_86_2_n_639 & csa_tree_add_86_2_n_630)));
 assign csa_tree_add_86_2_n_739 = (csa_tree_add_86_2_n_654 ^ (csa_tree_add_86_2_n_639 ^ csa_tree_add_86_2_n_630));
 assign csa_tree_add_86_2_n_736 = ((csa_tree_add_86_2_n_665 & csa_tree_add_86_2_n_632) | ((csa_tree_add_86_2_n_632
    & csa_tree_add_86_2_n_657) | (csa_tree_add_86_2_n_657 & csa_tree_add_86_2_n_665)));
 assign csa_tree_add_86_2_n_737 = (csa_tree_add_86_2_n_632 ^ (csa_tree_add_86_2_n_657 ^ csa_tree_add_86_2_n_665));
 assign csa_tree_add_86_2_n_734 = ((csa_tree_add_86_2_n_680 & csa_tree_add_86_2_n_603) | ((csa_tree_add_86_2_n_603
    & csa_tree_add_86_2_n_566) | (csa_tree_add_86_2_n_566 & csa_tree_add_86_2_n_680)));
 assign csa_tree_add_86_2_n_735 = (csa_tree_add_86_2_n_603 ^ (csa_tree_add_86_2_n_566 ^ csa_tree_add_86_2_n_680));
 assign csa_tree_add_86_2_n_732 = ((csa_tree_add_86_2_n_678 & csa_tree_add_86_2_n_567) | ((csa_tree_add_86_2_n_567
    & csa_tree_add_86_2_n_586) | (csa_tree_add_86_2_n_586 & csa_tree_add_86_2_n_678)));
 assign csa_tree_add_86_2_n_733 = (csa_tree_add_86_2_n_567 ^ (csa_tree_add_86_2_n_586 ^ csa_tree_add_86_2_n_678));
 assign csa_tree_add_86_2_n_730 = ((csa_tree_add_86_2_n_648 & csa_tree_add_86_2_n_620) | ((csa_tree_add_86_2_n_620
    & csa_tree_add_86_2_n_629) | (csa_tree_add_86_2_n_629 & csa_tree_add_86_2_n_648)));
 assign csa_tree_add_86_2_n_731 = (csa_tree_add_86_2_n_620 ^ (csa_tree_add_86_2_n_629 ^ csa_tree_add_86_2_n_648));
 assign csa_tree_add_86_2_n_728 = ((csa_tree_add_86_2_n_676 & csa_tree_add_86_2_n_590) | ((csa_tree_add_86_2_n_590
    & csa_tree_add_86_2_n_597) | (csa_tree_add_86_2_n_597 & csa_tree_add_86_2_n_676)));
 assign csa_tree_add_86_2_n_729 = (csa_tree_add_86_2_n_590 ^ (csa_tree_add_86_2_n_597 ^ csa_tree_add_86_2_n_676));
 assign csa_tree_add_86_2_n_726 = ((csa_tree_add_86_2_n_667 & csa_tree_add_86_2_n_623) | ((csa_tree_add_86_2_n_623
    & csa_tree_add_86_2_n_634) | (csa_tree_add_86_2_n_634 & csa_tree_add_86_2_n_667)));
 assign csa_tree_add_86_2_n_727 = (csa_tree_add_86_2_n_623 ^ (csa_tree_add_86_2_n_634 ^ csa_tree_add_86_2_n_667));
 assign csa_tree_add_86_2_n_724 = ((csa_tree_add_86_2_n_662 & csa_tree_add_86_2_n_658) | ((csa_tree_add_86_2_n_658
    & csa_tree_add_86_2_n_645) | (csa_tree_add_86_2_n_645 & csa_tree_add_86_2_n_662)));
 assign csa_tree_add_86_2_n_725 = (csa_tree_add_86_2_n_658 ^ (csa_tree_add_86_2_n_645 ^ csa_tree_add_86_2_n_662));
 assign csa_tree_add_86_2_n_722 = ((csa_tree_add_86_2_n_671 & csa_tree_add_86_2_n_485) | ((csa_tree_add_86_2_n_485
    & csa_tree_add_86_2_n_577) | (csa_tree_add_86_2_n_577 & csa_tree_add_86_2_n_671)));
 assign csa_tree_add_86_2_n_723 = (csa_tree_add_86_2_n_485 ^ (csa_tree_add_86_2_n_577 ^ csa_tree_add_86_2_n_671));
 assign csa_tree_add_86_2_n_720 = ((csa_tree_add_86_2_n_672 & csa_tree_add_86_2_n_581) | ((csa_tree_add_86_2_n_581
    & csa_tree_add_86_2_n_596) | (csa_tree_add_86_2_n_596 & csa_tree_add_86_2_n_672)));
 assign csa_tree_add_86_2_n_721 = (csa_tree_add_86_2_n_581 ^ (csa_tree_add_86_2_n_596 ^ csa_tree_add_86_2_n_672));
 assign csa_tree_add_86_2_n_718 = ((csa_tree_add_86_2_n_633 & csa_tree_add_86_2_n_227) | ((csa_tree_add_86_2_n_227
    & csa_tree_add_86_2_n_650) | (csa_tree_add_86_2_n_650 & csa_tree_add_86_2_n_633)));
 assign csa_tree_add_86_2_n_719 = (csa_tree_add_86_2_n_227 ^ (csa_tree_add_86_2_n_650 ^ csa_tree_add_86_2_n_633));
 assign csa_tree_add_86_2_n_716 = ((csa_tree_add_86_2_n_666 & csa_tree_add_86_2_n_587) | ((csa_tree_add_86_2_n_587
    & csa_tree_add_86_2_n_559) | (csa_tree_add_86_2_n_559 & csa_tree_add_86_2_n_666)));
 assign csa_tree_add_86_2_n_717 = (csa_tree_add_86_2_n_587 ^ (csa_tree_add_86_2_n_559 ^ csa_tree_add_86_2_n_666));
 assign csa_tree_add_86_2_n_714 = ((csa_tree_add_86_2_n_621 & csa_tree_add_86_2_n_589) | ((csa_tree_add_86_2_n_589
    & csa_tree_add_86_2_n_614) | (csa_tree_add_86_2_n_614 & csa_tree_add_86_2_n_621)));
 assign csa_tree_add_86_2_n_715 = (csa_tree_add_86_2_n_589 ^ (csa_tree_add_86_2_n_614 ^ csa_tree_add_86_2_n_621));
 assign csa_tree_add_86_2_n_712 = ((csa_tree_add_86_2_n_612 & csa_tree_add_86_2_n_617) | ((csa_tree_add_86_2_n_617
    & csa_tree_add_86_2_n_615) | (csa_tree_add_86_2_n_615 & csa_tree_add_86_2_n_612)));
 assign csa_tree_add_86_2_n_713 = (csa_tree_add_86_2_n_617 ^ (csa_tree_add_86_2_n_615 ^ csa_tree_add_86_2_n_612));
 assign csa_tree_add_86_2_n_710 = ((csa_tree_add_86_2_n_613 & csa_tree_add_86_2_n_95) | ((csa_tree_add_86_2_n_95
    & csa_tree_add_86_2_n_595) | (csa_tree_add_86_2_n_595 & csa_tree_add_86_2_n_613)));
 assign csa_tree_add_86_2_n_711 = (csa_tree_add_86_2_n_95 ^ (csa_tree_add_86_2_n_595 ^ csa_tree_add_86_2_n_613));
 assign csa_tree_add_86_2_n_708 = ((csa_tree_add_86_2_n_641 & csa_tree_add_86_2_n_579) | ((csa_tree_add_86_2_n_579
    & csa_tree_add_86_2_n_604) | (csa_tree_add_86_2_n_604 & csa_tree_add_86_2_n_641)));
 assign csa_tree_add_86_2_n_709 = (csa_tree_add_86_2_n_579 ^ (csa_tree_add_86_2_n_604 ^ csa_tree_add_86_2_n_641));
 assign csa_tree_add_86_2_n_706 = ((csa_tree_add_86_2_n_661 & csa_tree_add_86_2_n_184) | ((csa_tree_add_86_2_n_184
    & csa_tree_add_86_2_n_600) | (csa_tree_add_86_2_n_600 & csa_tree_add_86_2_n_661)));
 assign n_1405 = (csa_tree_add_86_2_n_184 ^ (csa_tree_add_86_2_n_600 ^ csa_tree_add_86_2_n_661));
 assign csa_tree_add_86_2_n_704 = ((csa_tree_add_86_2_n_619 & csa_tree_add_86_2_n_443) | ((csa_tree_add_86_2_n_443
    & csa_tree_add_86_2_n_580) | (csa_tree_add_86_2_n_580 & csa_tree_add_86_2_n_619)));
 assign csa_tree_add_86_2_n_705 = (csa_tree_add_86_2_n_443 ^ (csa_tree_add_86_2_n_580 ^ csa_tree_add_86_2_n_619));
 assign csa_tree_add_86_2_n_702 = ((csa_tree_add_86_2_n_610 & csa_tree_add_86_2_n_565) | ((csa_tree_add_86_2_n_565
    & csa_tree_add_86_2_n_509) | (csa_tree_add_86_2_n_509 & csa_tree_add_86_2_n_610)));
 assign csa_tree_add_86_2_n_703 = (csa_tree_add_86_2_n_565 ^ (csa_tree_add_86_2_n_509 ^ csa_tree_add_86_2_n_610));
 assign csa_tree_add_86_2_n_700 = ((csa_tree_add_86_2_n_592 & csa_tree_add_86_2_n_628) | ((csa_tree_add_86_2_n_628
    & csa_tree_add_86_2_n_514) | (csa_tree_add_86_2_n_514 & csa_tree_add_86_2_n_592)));
 assign csa_tree_add_86_2_n_701 = (csa_tree_add_86_2_n_628 ^ (csa_tree_add_86_2_n_514 ^ csa_tree_add_86_2_n_592));
 assign csa_tree_add_86_2_n_698 = ((csa_tree_add_86_2_n_644 & csa_tree_add_86_2_n_506) | ((csa_tree_add_86_2_n_506
    & csa_tree_add_86_2_n_521) | (csa_tree_add_86_2_n_521 & csa_tree_add_86_2_n_644)));
 assign csa_tree_add_86_2_n_699 = (csa_tree_add_86_2_n_506 ^ (csa_tree_add_86_2_n_521 ^ csa_tree_add_86_2_n_644));
 assign csa_tree_add_86_2_n_696 = ((csa_tree_add_86_2_n_616 & csa_tree_add_86_2_n_523) | ((csa_tree_add_86_2_n_523
    & csa_tree_add_86_2_n_582) | (csa_tree_add_86_2_n_582 & csa_tree_add_86_2_n_616)));
 assign csa_tree_add_86_2_n_697 = (csa_tree_add_86_2_n_523 ^ (csa_tree_add_86_2_n_582 ^ csa_tree_add_86_2_n_616));
 assign csa_tree_add_86_2_n_694 = ((csa_tree_add_86_2_n_627 & csa_tree_add_86_2_n_126) | ((csa_tree_add_86_2_n_126
    & csa_tree_add_86_2_n_593) | (csa_tree_add_86_2_n_593 & csa_tree_add_86_2_n_627)));
 assign csa_tree_add_86_2_n_695 = (csa_tree_add_86_2_n_126 ^ (csa_tree_add_86_2_n_593 ^ csa_tree_add_86_2_n_627));
 assign csa_tree_add_86_2_n_692 = ((csa_tree_add_86_2_n_642 & csa_tree_add_86_2_n_584) | ((csa_tree_add_86_2_n_584
    & csa_tree_add_86_2_n_591) | (csa_tree_add_86_2_n_591 & csa_tree_add_86_2_n_642)));
 assign csa_tree_add_86_2_n_693 = (csa_tree_add_86_2_n_584 ^ (csa_tree_add_86_2_n_591 ^ csa_tree_add_86_2_n_642));
 assign csa_tree_add_86_2_n_690 = ((csa_tree_add_86_2_n_640 & csa_tree_add_86_2_n_578) | ((csa_tree_add_86_2_n_578
    & csa_tree_add_86_2_n_483) | (csa_tree_add_86_2_n_483 & csa_tree_add_86_2_n_640)));
 assign csa_tree_add_86_2_n_691 = (csa_tree_add_86_2_n_578 ^ (csa_tree_add_86_2_n_483 ^ csa_tree_add_86_2_n_640));
 assign csa_tree_add_86_2_n_688 = ((csa_tree_add_86_2_n_576 & csa_tree_add_86_2_n_484) | ((csa_tree_add_86_2_n_484
    & csa_tree_add_86_2_n_553) | (csa_tree_add_86_2_n_553 & csa_tree_add_86_2_n_576)));
 assign csa_tree_add_86_2_n_689 = (csa_tree_add_86_2_n_484 ^ (csa_tree_add_86_2_n_553 ^ csa_tree_add_86_2_n_576));
 assign csa_tree_add_86_2_n_686 = ((csa_tree_add_86_2_n_598 & csa_tree_add_86_2_n_451) | ((csa_tree_add_86_2_n_451
    & csa_tree_add_86_2_n_519) | (csa_tree_add_86_2_n_519 & csa_tree_add_86_2_n_598)));
 assign csa_tree_add_86_2_n_687 = (csa_tree_add_86_2_n_451 ^ (csa_tree_add_86_2_n_519 ^ csa_tree_add_86_2_n_598));
 assign csa_tree_add_86_2_n_684 = ((csa_tree_add_86_2_n_575 & csa_tree_add_86_2_n_564) | ((csa_tree_add_86_2_n_564
    & csa_tree_add_86_2_n_481) | (csa_tree_add_86_2_n_481 & csa_tree_add_86_2_n_575)));
 assign csa_tree_add_86_2_n_685 = (csa_tree_add_86_2_n_564 ^ (csa_tree_add_86_2_n_481 ^ csa_tree_add_86_2_n_575));
 assign csa_tree_add_86_2_n_682 = ((csa_tree_add_86_2_n_618 & csa_tree_add_86_2_n_448) | ((csa_tree_add_86_2_n_448
    & csa_tree_add_86_2_n_461) | (csa_tree_add_86_2_n_461 & csa_tree_add_86_2_n_618)));
 assign csa_tree_add_86_2_n_683 = (csa_tree_add_86_2_n_448 ^ (csa_tree_add_86_2_n_461 ^ csa_tree_add_86_2_n_618));
 assign csa_tree_add_86_2_n_680 = ((csa_tree_add_86_2_n_599 & csa_tree_add_86_2_n_558) | ((csa_tree_add_86_2_n_558
    & csa_tree_add_86_2_n_471) | (csa_tree_add_86_2_n_471 & csa_tree_add_86_2_n_599)));
 assign csa_tree_add_86_2_n_681 = (csa_tree_add_86_2_n_558 ^ (csa_tree_add_86_2_n_471 ^ csa_tree_add_86_2_n_599));
 assign csa_tree_add_86_2_n_678 = ((csa_tree_add_86_2_n_622 & csa_tree_add_86_2_n_446) | ((csa_tree_add_86_2_n_446
    & csa_tree_add_86_2_n_455) | (csa_tree_add_86_2_n_455 & csa_tree_add_86_2_n_622)));
 assign csa_tree_add_86_2_n_679 = (csa_tree_add_86_2_n_446 ^ (csa_tree_add_86_2_n_455 ^ csa_tree_add_86_2_n_622));
 assign csa_tree_add_86_2_n_676 = ((csa_tree_add_86_2_n_573 & csa_tree_add_86_2_n_562) | ((csa_tree_add_86_2_n_562
    & csa_tree_add_86_2_n_429) | (csa_tree_add_86_2_n_429 & csa_tree_add_86_2_n_573)));
 assign csa_tree_add_86_2_n_677 = (csa_tree_add_86_2_n_562 ^ (csa_tree_add_86_2_n_429 ^ csa_tree_add_86_2_n_573));
 assign csa_tree_add_86_2_n_674 = ((csa_tree_add_86_2_n_583 & csa_tree_add_86_2_n_594) | ((csa_tree_add_86_2_n_594
    & csa_tree_add_86_2_n_482) | (csa_tree_add_86_2_n_482 & csa_tree_add_86_2_n_583)));
 assign csa_tree_add_86_2_n_675 = (csa_tree_add_86_2_n_594 ^ (csa_tree_add_86_2_n_482 ^ csa_tree_add_86_2_n_583));
 assign csa_tree_add_86_2_n_672 = ((csa_tree_add_86_2_n_457 & csa_tree_add_86_2_n_445) | ((csa_tree_add_86_2_n_445
    & csa_tree_add_86_2_n_572) | (csa_tree_add_86_2_n_572 & csa_tree_add_86_2_n_457)));
 assign csa_tree_add_86_2_n_673 = (csa_tree_add_86_2_n_445 ^ (csa_tree_add_86_2_n_572 ^ csa_tree_add_86_2_n_457));
 assign csa_tree_add_86_2_n_670 = ((csa_tree_add_86_2_n_571 & csa_tree_add_86_2_n_606) | ((csa_tree_add_86_2_n_606
    & csa_tree_add_86_2_n_574) | (csa_tree_add_86_2_n_574 & csa_tree_add_86_2_n_571)));
 assign csa_tree_add_86_2_n_671 = (csa_tree_add_86_2_n_606 ^ (csa_tree_add_86_2_n_574 ^ csa_tree_add_86_2_n_571));
 assign csa_tree_add_86_2_n_666 = ((csa_tree_add_86_2_n_560 & csa_tree_add_86_2_n_447) | ((csa_tree_add_86_2_n_447
    & csa_tree_add_86_2_n_503) | (csa_tree_add_86_2_n_503 & csa_tree_add_86_2_n_560)));
 assign csa_tree_add_86_2_n_667 = (csa_tree_add_86_2_n_447 ^ (csa_tree_add_86_2_n_503 ^ csa_tree_add_86_2_n_560));
 assign csa_tree_add_86_2_n_664 = ((csa_tree_add_86_2_n_513 & csa_tree_add_86_2_n_458) | ((csa_tree_add_86_2_n_458
    & csa_tree_add_86_2_n_541) | (csa_tree_add_86_2_n_541 & csa_tree_add_86_2_n_513)));
 assign csa_tree_add_86_2_n_665 = (csa_tree_add_86_2_n_458 ^ (csa_tree_add_86_2_n_541 ^ csa_tree_add_86_2_n_513));
 assign csa_tree_add_86_2_n_662 = ((csa_tree_add_86_2_n_505 & csa_tree_add_86_2_n_530) | ((csa_tree_add_86_2_n_530
    & csa_tree_add_86_2_n_501) | (csa_tree_add_86_2_n_501 & csa_tree_add_86_2_n_505)));
 assign csa_tree_add_86_2_n_663 = (csa_tree_add_86_2_n_530 ^ (csa_tree_add_86_2_n_501 ^ csa_tree_add_86_2_n_505));
 assign csa_tree_add_86_2_n_660 = ((csa_tree_add_86_2_n_605 & csa_tree_add_86_2_n_516) | ((csa_tree_add_86_2_n_516
    & csa_tree_add_86_2_n_479) | (csa_tree_add_86_2_n_479 & csa_tree_add_86_2_n_605)));
 assign csa_tree_add_86_2_n_661 = (csa_tree_add_86_2_n_516 ^ (csa_tree_add_86_2_n_479 ^ csa_tree_add_86_2_n_605));
 assign csa_tree_add_86_2_n_658 = ((csa_tree_add_86_2_n_512 & csa_tree_add_86_2_n_540) | ((csa_tree_add_86_2_n_540
    & csa_tree_add_86_2_n_536) | (csa_tree_add_86_2_n_536 & csa_tree_add_86_2_n_512)));
 assign csa_tree_add_86_2_n_659 = (csa_tree_add_86_2_n_540 ^ (csa_tree_add_86_2_n_536 ^ csa_tree_add_86_2_n_512));
 assign csa_tree_add_86_2_n_656 = ((csa_tree_add_86_2_n_534 & csa_tree_add_86_2_n_531) | ((csa_tree_add_86_2_n_531
    & csa_tree_add_86_2_n_537) | (csa_tree_add_86_2_n_537 & csa_tree_add_86_2_n_534)));
 assign csa_tree_add_86_2_n_657 = (csa_tree_add_86_2_n_531 ^ (csa_tree_add_86_2_n_537 ^ csa_tree_add_86_2_n_534));
 assign csa_tree_add_86_2_n_654 = ((csa_tree_add_86_2_n_494 & csa_tree_add_86_2_n_538) | ((csa_tree_add_86_2_n_538
    & csa_tree_add_86_2_n_532) | (csa_tree_add_86_2_n_532 & csa_tree_add_86_2_n_494)));
 assign csa_tree_add_86_2_n_655 = (csa_tree_add_86_2_n_538 ^ (csa_tree_add_86_2_n_532 ^ csa_tree_add_86_2_n_494));
 assign csa_tree_add_86_2_n_652 = ((csa_tree_add_86_2_n_492 & csa_tree_add_86_2_n_263) | ((csa_tree_add_86_2_n_263
    & csa_tree_add_86_2_n_520) | (csa_tree_add_86_2_n_520 & csa_tree_add_86_2_n_492)));
 assign csa_tree_add_86_2_n_653 = (csa_tree_add_86_2_n_263 ^ (csa_tree_add_86_2_n_520 ^ csa_tree_add_86_2_n_492));
 assign csa_tree_add_86_2_n_650 = ((csa_tree_add_86_2_n_588 & csa_tree_add_86_2_n_539) | ((csa_tree_add_86_2_n_539
    & csa_tree_add_86_2_n_515) | (csa_tree_add_86_2_n_515 & csa_tree_add_86_2_n_588)));
 assign csa_tree_add_86_2_n_651 = (csa_tree_add_86_2_n_539 ^ (csa_tree_add_86_2_n_515 ^ csa_tree_add_86_2_n_588));
 assign csa_tree_add_86_2_n_648 = ((csa_tree_add_86_2_n_499 & csa_tree_add_86_2_n_543) | ((csa_tree_add_86_2_n_543
    & csa_tree_add_86_2_n_489) | (csa_tree_add_86_2_n_489 & csa_tree_add_86_2_n_499)));
 assign csa_tree_add_86_2_n_649 = (csa_tree_add_86_2_n_543 ^ (csa_tree_add_86_2_n_489 ^ csa_tree_add_86_2_n_499));
 assign csa_tree_add_86_2_n_646 = ((csa_tree_add_86_2_n_507 & csa_tree_add_86_2_n_524) | ((csa_tree_add_86_2_n_524
    & csa_tree_add_86_2_n_477) | (csa_tree_add_86_2_n_477 & csa_tree_add_86_2_n_507)));
 assign csa_tree_add_86_2_n_647 = (csa_tree_add_86_2_n_524 ^ (csa_tree_add_86_2_n_477 ^ csa_tree_add_86_2_n_507));
 assign csa_tree_add_86_2_n_644 = ((csa_tree_add_86_2_n_475 & csa_tree_add_86_2_n_504) | ((csa_tree_add_86_2_n_504
    & csa_tree_add_86_2_n_500) | (csa_tree_add_86_2_n_500 & csa_tree_add_86_2_n_475)));
 assign csa_tree_add_86_2_n_645 = (csa_tree_add_86_2_n_504 ^ (csa_tree_add_86_2_n_500 ^ csa_tree_add_86_2_n_475));
 assign csa_tree_add_86_2_n_642 = ((csa_tree_add_86_2_n_563 & csa_tree_add_86_2_n_518) | ((csa_tree_add_86_2_n_518
    & csa_tree_add_86_2_n_439) | (csa_tree_add_86_2_n_439 & csa_tree_add_86_2_n_563)));
 assign csa_tree_add_86_2_n_643 = (csa_tree_add_86_2_n_518 ^ (csa_tree_add_86_2_n_439 ^ csa_tree_add_86_2_n_563));
 assign csa_tree_add_86_2_n_640 = ((csa_tree_add_86_2_n_491 & csa_tree_add_86_2_n_545) | ((csa_tree_add_86_2_n_545
    & csa_tree_add_86_2_n_478) | (csa_tree_add_86_2_n_478 & csa_tree_add_86_2_n_491)));
 assign csa_tree_add_86_2_n_641 = (csa_tree_add_86_2_n_545 ^ (csa_tree_add_86_2_n_478 ^ csa_tree_add_86_2_n_491));
 assign csa_tree_add_86_2_n_638 = ((csa_tree_add_86_2_n_472 & csa_tree_add_86_2_n_430) | ((csa_tree_add_86_2_n_430
    & csa_tree_add_86_2_n_468) | (csa_tree_add_86_2_n_468 & csa_tree_add_86_2_n_472)));
 assign csa_tree_add_86_2_n_639 = (csa_tree_add_86_2_n_430 ^ (csa_tree_add_86_2_n_468 ^ csa_tree_add_86_2_n_472));
 assign csa_tree_add_86_2_n_636 = ((csa_tree_add_86_2_n_453 & csa_tree_add_86_2_n_444) | ((csa_tree_add_86_2_n_444
    & csa_tree_add_86_2_n_435) | (csa_tree_add_86_2_n_435 & csa_tree_add_86_2_n_453)));
 assign csa_tree_add_86_2_n_637 = (csa_tree_add_86_2_n_444 ^ (csa_tree_add_86_2_n_435 ^ csa_tree_add_86_2_n_453));
 assign csa_tree_add_86_2_n_634 = ((csa_tree_add_86_2_n_570 & csa_tree_add_86_2_n_187) | ((csa_tree_add_86_2_n_187
    & csa_tree_add_86_2_n_185) | (csa_tree_add_86_2_n_185 & csa_tree_add_86_2_n_570)));
 assign csa_tree_add_86_2_n_635 = (csa_tree_add_86_2_n_187 ^ (csa_tree_add_86_2_n_185 ^ csa_tree_add_86_2_n_570));
 assign csa_tree_add_86_2_n_632 = ((csa_tree_add_86_2_n_535 & csa_tree_add_86_2_n_473) | ((csa_tree_add_86_2_n_473
    & csa_tree_add_86_2_n_431) | (csa_tree_add_86_2_n_431 & csa_tree_add_86_2_n_535)));
 assign csa_tree_add_86_2_n_633 = (csa_tree_add_86_2_n_473 ^ (csa_tree_add_86_2_n_431 ^ csa_tree_add_86_2_n_535));
 assign csa_tree_add_86_2_n_630 = ((csa_tree_add_86_2_n_469 & csa_tree_add_86_2_n_528) | ((csa_tree_add_86_2_n_528
    & csa_tree_add_86_2_n_459) | (csa_tree_add_86_2_n_459 & csa_tree_add_86_2_n_469)));
 assign csa_tree_add_86_2_n_631 = (csa_tree_add_86_2_n_528 ^ (csa_tree_add_86_2_n_459 ^ csa_tree_add_86_2_n_469));
 assign csa_tree_add_86_2_n_628 = ((csa_tree_add_86_2_n_522 & csa_tree_add_86_2_n_498) | ((csa_tree_add_86_2_n_498
    & csa_tree_add_86_2_n_542) | (csa_tree_add_86_2_n_542 & csa_tree_add_86_2_n_522)));
 assign csa_tree_add_86_2_n_629 = (csa_tree_add_86_2_n_498 ^ (csa_tree_add_86_2_n_542 ^ csa_tree_add_86_2_n_522));
 assign csa_tree_add_86_2_n_626 = ((csa_tree_add_86_2_n_529 & csa_tree_add_86_2_n_533) | ((csa_tree_add_86_2_n_533
    & csa_tree_add_86_2_n_495) | (csa_tree_add_86_2_n_495 & csa_tree_add_86_2_n_529)));
 assign csa_tree_add_86_2_n_627 = (csa_tree_add_86_2_n_533 ^ (csa_tree_add_86_2_n_495 ^ csa_tree_add_86_2_n_529));
 assign csa_tree_add_86_2_n_624 = ((csa_tree_add_86_2_n_493 & csa_tree_add_86_2_n_474) | ((csa_tree_add_86_2_n_474
    & csa_tree_add_86_2_n_476) | (csa_tree_add_86_2_n_476 & csa_tree_add_86_2_n_493)));
 assign csa_tree_add_86_2_n_625 = (csa_tree_add_86_2_n_474 ^ (csa_tree_add_86_2_n_476 ^ csa_tree_add_86_2_n_493));
 assign csa_tree_add_86_2_n_622 = ((csa_tree_add_86_2_n_552 & csa_tree_add_86_2_n_170) | ((csa_tree_add_86_2_n_170
    & csa_tree_add_86_2_n_417) | (csa_tree_add_86_2_n_417 & csa_tree_add_86_2_n_552)));
 assign csa_tree_add_86_2_n_623 = (csa_tree_add_86_2_n_170 ^ (csa_tree_add_86_2_n_417 ^ csa_tree_add_86_2_n_552));
 assign csa_tree_add_86_2_n_620 = ((csa_tree_add_86_2_n_486 & csa_tree_add_86_2_n_223) | ((csa_tree_add_86_2_n_223
    & csa_tree_add_86_2_n_510) | (csa_tree_add_86_2_n_510 & csa_tree_add_86_2_n_486)));
 assign csa_tree_add_86_2_n_621 = (csa_tree_add_86_2_n_223 ^ (csa_tree_add_86_2_n_510 ^ csa_tree_add_86_2_n_486));
 assign csa_tree_add_86_2_n_618 = ((csa_tree_add_86_2_n_449 & csa_tree_add_86_2_n_452) | ((csa_tree_add_86_2_n_452
    & csa_tree_add_86_2_n_434) | (csa_tree_add_86_2_n_434 & csa_tree_add_86_2_n_449)));
 assign csa_tree_add_86_2_n_619 = (csa_tree_add_86_2_n_452 ^ (csa_tree_add_86_2_n_434 ^ csa_tree_add_86_2_n_449));
 assign csa_tree_add_86_2_n_616 = ((csa_tree_add_86_2_n_546 & csa_tree_add_86_2_n_91) | ((csa_tree_add_86_2_n_91
    & csa_tree_add_86_2_n_496) | (csa_tree_add_86_2_n_496 & csa_tree_add_86_2_n_546)));
 assign csa_tree_add_86_2_n_617 = (csa_tree_add_86_2_n_91 ^ (csa_tree_add_86_2_n_496 ^ csa_tree_add_86_2_n_546));
 assign csa_tree_add_86_2_n_614 = ((csa_tree_add_86_2_n_527 & csa_tree_add_86_2_n_487) | ((csa_tree_add_86_2_n_487
    & csa_tree_add_86_2_n_511) | (csa_tree_add_86_2_n_511 & csa_tree_add_86_2_n_527)));
 assign csa_tree_add_86_2_n_615 = (csa_tree_add_86_2_n_487 ^ (csa_tree_add_86_2_n_511 ^ csa_tree_add_86_2_n_527));
 assign csa_tree_add_86_2_n_612 = ((csa_tree_add_86_2_n_497 & csa_tree_add_86_2_n_544) | ((csa_tree_add_86_2_n_544
    & csa_tree_add_86_2_n_547) | (csa_tree_add_86_2_n_547 & csa_tree_add_86_2_n_497)));
 assign csa_tree_add_86_2_n_613 = (csa_tree_add_86_2_n_544 ^ (csa_tree_add_86_2_n_547 ^ csa_tree_add_86_2_n_497));
 assign csa_tree_add_86_2_n_610 = ((csa_tree_add_86_2_n_391 & csa_tree_add_86_2_n_137) | ((csa_tree_add_86_2_n_137
    & csa_tree_add_86_2_n_440) | (csa_tree_add_86_2_n_440 & csa_tree_add_86_2_n_391)));
 assign csa_tree_add_86_2_n_611 = (csa_tree_add_86_2_n_137 ^ (csa_tree_add_86_2_n_440 ^ csa_tree_add_86_2_n_391));
 assign csa_tree_add_86_2_n_606 = ((csa_tree_add_86_2_n_508 & csa_tree_add_86_2_n_63) | ((csa_tree_add_86_2_n_63
    & csa_tree_add_86_2_n_96) | (csa_tree_add_86_2_n_96 & csa_tree_add_86_2_n_508)));
 assign csa_tree_add_86_2_n_607 = (csa_tree_add_86_2_n_63 ^ (csa_tree_add_86_2_n_96 ^ csa_tree_add_86_2_n_508));
 assign csa_tree_add_86_2_n_604 = ((csa_tree_add_86_2_n_549 & csa_tree_add_86_2_n_84) | ((csa_tree_add_86_2_n_84
    & csa_tree_add_86_2_n_404) | (csa_tree_add_86_2_n_404 & csa_tree_add_86_2_n_549)));
 assign csa_tree_add_86_2_n_605 = (csa_tree_add_86_2_n_84 ^ (csa_tree_add_86_2_n_404 ^ csa_tree_add_86_2_n_549));
 assign csa_tree_add_86_2_n_602 = ((csa_tree_add_86_2_n_470 & csa_tree_add_86_2_n_149) | ((csa_tree_add_86_2_n_149
    & csa_tree_add_86_2_n_395) | (csa_tree_add_86_2_n_395 & csa_tree_add_86_2_n_470)));
 assign csa_tree_add_86_2_n_603 = (csa_tree_add_86_2_n_149 ^ (csa_tree_add_86_2_n_395 ^ csa_tree_add_86_2_n_470));
 assign csa_tree_add_86_2_n_600 = ((csa_tree_add_86_2_n_517 & csa_tree_add_86_2_n_72) | ((csa_tree_add_86_2_n_72
    & csa_tree_add_86_2_n_405) | (csa_tree_add_86_2_n_405 & csa_tree_add_86_2_n_517)));
 assign n_1406 = (csa_tree_add_86_2_n_72 ^ (csa_tree_add_86_2_n_405 ^ csa_tree_add_86_2_n_517));
 assign csa_tree_add_86_2_n_598 = ((csa_tree_add_86_2_n_413 & csa_tree_add_86_2_n_97) | ((csa_tree_add_86_2_n_97
    & csa_tree_add_86_2_n_408) | (csa_tree_add_86_2_n_408 & csa_tree_add_86_2_n_413)));
 assign csa_tree_add_86_2_n_599 = (csa_tree_add_86_2_n_97 ^ (csa_tree_add_86_2_n_408 ^ csa_tree_add_86_2_n_413));
 assign csa_tree_add_86_2_n_596 = ((csa_tree_add_86_2_n_428 & csa_tree_add_86_2_n_415) | ((csa_tree_add_86_2_n_415
    & csa_tree_add_86_2_n_422) | (csa_tree_add_86_2_n_422 & csa_tree_add_86_2_n_428)));
 assign csa_tree_add_86_2_n_597 = (csa_tree_add_86_2_n_415 ^ (csa_tree_add_86_2_n_422 ^ csa_tree_add_86_2_n_428));
 assign csa_tree_add_86_2_n_594 = ((csa_tree_add_86_2_n_490 & csa_tree_add_86_2_n_189) | ((csa_tree_add_86_2_n_189
    & csa_tree_add_86_2_n_425) | (csa_tree_add_86_2_n_425 & csa_tree_add_86_2_n_490)));
 assign csa_tree_add_86_2_n_595 = (csa_tree_add_86_2_n_189 ^ (csa_tree_add_86_2_n_425 ^ csa_tree_add_86_2_n_490));
 assign csa_tree_add_86_2_n_592 = ((csa_tree_add_86_2_n_488 & csa_tree_add_86_2_n_249) | ((csa_tree_add_86_2_n_249
    & csa_tree_add_86_2_n_420) | (csa_tree_add_86_2_n_420 & csa_tree_add_86_2_n_488)));
 assign csa_tree_add_86_2_n_593 = (csa_tree_add_86_2_n_249 ^ (csa_tree_add_86_2_n_420 ^ csa_tree_add_86_2_n_488));
 assign csa_tree_add_86_2_n_590 = ((csa_tree_add_86_2_n_438 & csa_tree_add_86_2_n_298) | ((csa_tree_add_86_2_n_298
    & csa_tree_add_86_2_n_423) | (csa_tree_add_86_2_n_423 & csa_tree_add_86_2_n_438)));
 assign csa_tree_add_86_2_n_591 = (csa_tree_add_86_2_n_298 ^ (csa_tree_add_86_2_n_423 ^ csa_tree_add_86_2_n_438));
 assign csa_tree_add_86_2_n_588 = ((csa_tree_add_86_2_n_526 & csa_tree_add_86_2_n_418) | ((csa_tree_add_86_2_n_418
    & csa_tree_add_86_2_n_421) | (csa_tree_add_86_2_n_421 & csa_tree_add_86_2_n_526)));
 assign csa_tree_add_86_2_n_589 = (csa_tree_add_86_2_n_418 ^ (csa_tree_add_86_2_n_421 ^ csa_tree_add_86_2_n_526));
 assign csa_tree_add_86_2_n_586 = ((csa_tree_add_86_2_n_502 & csa_tree_add_86_2_n_180) | ((csa_tree_add_86_2_n_180
    & csa_tree_add_86_2_n_39) | (csa_tree_add_86_2_n_39 & csa_tree_add_86_2_n_502)));
 assign csa_tree_add_86_2_n_587 = (csa_tree_add_86_2_n_180 ^ (csa_tree_add_86_2_n_39 ^ csa_tree_add_86_2_n_502));
 assign csa_tree_add_86_2_n_584 = ((csa_tree_add_86_2_n_450 & csa_tree_add_86_2_n_112) | ((csa_tree_add_86_2_n_112
    & csa_tree_add_86_2_n_394) | (csa_tree_add_86_2_n_394 & csa_tree_add_86_2_n_450)));
 assign csa_tree_add_86_2_n_585 = (csa_tree_add_86_2_n_112 ^ (csa_tree_add_86_2_n_394 ^ csa_tree_add_86_2_n_450));
 assign csa_tree_add_86_2_n_582 = ((csa_tree_add_86_2_n_419 & csa_tree_add_86_2_n_303) | ((csa_tree_add_86_2_n_303
    & csa_tree_add_86_2_n_424) | (csa_tree_add_86_2_n_424 & csa_tree_add_86_2_n_419)));
 assign csa_tree_add_86_2_n_583 = (csa_tree_add_86_2_n_303 ^ (csa_tree_add_86_2_n_424 ^ csa_tree_add_86_2_n_419));
 assign csa_tree_add_86_2_n_580 = ((csa_tree_add_86_2_n_456 & csa_tree_add_86_2_n_295) | ((csa_tree_add_86_2_n_295
    & csa_tree_add_86_2_n_414) | (csa_tree_add_86_2_n_414 & csa_tree_add_86_2_n_456)));
 assign csa_tree_add_86_2_n_581 = (csa_tree_add_86_2_n_295 ^ (csa_tree_add_86_2_n_414 ^ csa_tree_add_86_2_n_456));
 assign csa_tree_add_86_2_n_578 = ((csa_tree_add_86_2_n_548 & csa_tree_add_86_2_n_171) | ((csa_tree_add_86_2_n_171
    & csa_tree_add_86_2_n_403) | (csa_tree_add_86_2_n_403 & csa_tree_add_86_2_n_548)));
 assign csa_tree_add_86_2_n_579 = (csa_tree_add_86_2_n_171 ^ (csa_tree_add_86_2_n_403 ^ csa_tree_add_86_2_n_548));
 assign csa_tree_add_86_2_n_576 = ((csa_tree_add_86_2_n_480 & csa_tree_add_86_2_n_46) | ((csa_tree_add_86_2_n_46
    & csa_tree_add_86_2_n_50) | (csa_tree_add_86_2_n_50 & csa_tree_add_86_2_n_480)));
 assign csa_tree_add_86_2_n_577 = (csa_tree_add_86_2_n_46 ^ (csa_tree_add_86_2_n_50 ^ csa_tree_add_86_2_n_480));
 assign csa_tree_add_86_2_n_574 = ((csa_tree_add_86_2_n_389 & csa_tree_add_86_2_n_89) | ((csa_tree_add_86_2_n_89
    & csa_tree_add_86_2_n_80) | (csa_tree_add_86_2_n_80 & csa_tree_add_86_2_n_389)));
 assign csa_tree_add_86_2_n_575 = (csa_tree_add_86_2_n_89 ^ (csa_tree_add_86_2_n_80 ^ csa_tree_add_86_2_n_389));
 assign csa_tree_add_86_2_n_572 = ((csa_tree_add_86_2_n_406 & csa_tree_add_86_2_n_123) | ((csa_tree_add_86_2_n_123
    & csa_tree_add_86_2_n_155) | (csa_tree_add_86_2_n_155 & csa_tree_add_86_2_n_406)));
 assign csa_tree_add_86_2_n_573 = (csa_tree_add_86_2_n_123 ^ (csa_tree_add_86_2_n_155 ^ csa_tree_add_86_2_n_406));
 assign csa_tree_add_86_2_n_570 = ((csa_tree_add_86_2_n_388 & csa_tree_add_86_2_n_62) | ((csa_tree_add_86_2_n_62
    & csa_tree_add_86_2_n_128) | (csa_tree_add_86_2_n_128 & csa_tree_add_86_2_n_388)));
 assign csa_tree_add_86_2_n_571 = (csa_tree_add_86_2_n_62 ^ (csa_tree_add_86_2_n_128 ^ csa_tree_add_86_2_n_388));
 assign csa_tree_add_86_2_n_566 = ((csa_tree_add_86_2_n_454 & csa_tree_add_86_2_n_71) | ((csa_tree_add_86_2_n_71
    & csa_tree_add_86_2_n_45) | (csa_tree_add_86_2_n_45 & csa_tree_add_86_2_n_454)));
 assign csa_tree_add_86_2_n_567 = (csa_tree_add_86_2_n_71 ^ (csa_tree_add_86_2_n_45 ^ csa_tree_add_86_2_n_454));
 assign csa_tree_add_86_2_n_564 = ((csa_tree_add_86_2_n_393 & csa_tree_add_86_2_n_92) | ((csa_tree_add_86_2_n_92
    & csa_tree_add_86_2_n_129) | (csa_tree_add_86_2_n_129 & csa_tree_add_86_2_n_393)));
 assign csa_tree_add_86_2_n_565 = (csa_tree_add_86_2_n_92 ^ (csa_tree_add_86_2_n_129 ^ csa_tree_add_86_2_n_393));
 assign csa_tree_add_86_2_n_562 = ((csa_tree_add_86_2_n_407 & csa_tree_add_86_2_n_120) | ((csa_tree_add_86_2_n_120
    & csa_tree_add_86_2_n_176) | (csa_tree_add_86_2_n_176 & csa_tree_add_86_2_n_407)));
 assign csa_tree_add_86_2_n_563 = (csa_tree_add_86_2_n_120 ^ (csa_tree_add_86_2_n_176 ^ csa_tree_add_86_2_n_407));
 assign csa_tree_add_86_2_n_560 = ((csa_tree_add_86_2_n_427 & csa_tree_add_86_2_n_48) | ((csa_tree_add_86_2_n_48
    & csa_tree_add_86_2_n_168) | (csa_tree_add_86_2_n_168 & csa_tree_add_86_2_n_427)));
 assign csa_tree_add_86_2_n_561 = (csa_tree_add_86_2_n_48 ^ (csa_tree_add_86_2_n_168 ^ csa_tree_add_86_2_n_427));
 assign csa_tree_add_86_2_n_558 = ((csa_tree_add_86_2_n_416 & csa_tree_add_86_2_n_53) | ((csa_tree_add_86_2_n_53
    & csa_tree_add_86_2_n_409) | (csa_tree_add_86_2_n_409 & csa_tree_add_86_2_n_416)));
 assign csa_tree_add_86_2_n_559 = (csa_tree_add_86_2_n_53 ^ (csa_tree_add_86_2_n_409 ^ csa_tree_add_86_2_n_416));
 assign csa_tree_add_86_2_n_556 = ((csa_tree_add_86_2_n_466 & csa_tree_add_86_2_n_218) | ((csa_tree_add_86_2_n_218
    & csa_tree_add_86_2_n_256) | (csa_tree_add_86_2_n_256 & csa_tree_add_86_2_n_466)));
 assign csa_tree_add_86_2_n_557 = (csa_tree_add_86_2_n_218 ^ (csa_tree_add_86_2_n_256 ^ csa_tree_add_86_2_n_466));
 assign csa_tree_add_86_2_n_554 = ((csa_tree_add_86_2_n_442 & csa_tree_add_86_2_n_136) | ((csa_tree_add_86_2_n_136
    & csa_tree_add_86_2_n_277) | (csa_tree_add_86_2_n_277 & csa_tree_add_86_2_n_442)));
 assign csa_tree_add_86_2_n_555 = (csa_tree_add_86_2_n_136 ^ (csa_tree_add_86_2_n_277 ^ csa_tree_add_86_2_n_442));
 assign csa_tree_add_86_2_n_552 = ((csa_tree_add_86_2_n_410 & csa_tree_add_86_2_n_93) | ((csa_tree_add_86_2_n_93
    & csa_tree_add_86_2_n_78) | (csa_tree_add_86_2_n_78 & csa_tree_add_86_2_n_410)));
 assign csa_tree_add_86_2_n_553 = (csa_tree_add_86_2_n_93 ^ (csa_tree_add_86_2_n_78 ^ csa_tree_add_86_2_n_410));
 assign csa_tree_add_86_2_n_550 = ((csa_tree_add_86_2_n_462 & csa_tree_add_86_2_n_49) | ((csa_tree_add_86_2_n_49
    & csa_tree_add_86_2_n_102) | (csa_tree_add_86_2_n_102 & csa_tree_add_86_2_n_462)));
 assign csa_tree_add_86_2_n_551 = (csa_tree_add_86_2_n_49 ^ (csa_tree_add_86_2_n_102 ^ csa_tree_add_86_2_n_462));
 assign csa_tree_add_86_2_n_548 = ((csa_tree_add_86_2_n_350 & csa_tree_add_86_2_n_261) | ((csa_tree_add_86_2_n_261
    & csa_tree_add_86_2_n_262) | (csa_tree_add_86_2_n_262 & csa_tree_add_86_2_n_350)));
 assign csa_tree_add_86_2_n_549 = (csa_tree_add_86_2_n_261 ^ (csa_tree_add_86_2_n_262 ^ csa_tree_add_86_2_n_350));
 assign csa_tree_add_86_2_n_546 = ((csa_tree_add_86_2_n_345 & csa_tree_add_86_2_n_278) | ((csa_tree_add_86_2_n_278
    & csa_tree_add_86_2_n_257) | (csa_tree_add_86_2_n_257 & csa_tree_add_86_2_n_345)));
 assign csa_tree_add_86_2_n_547 = (csa_tree_add_86_2_n_278 ^ (csa_tree_add_86_2_n_257 ^ csa_tree_add_86_2_n_345));
 assign csa_tree_add_86_2_n_544 = ((csa_tree_add_86_2_n_327 & csa_tree_add_86_2_n_269) | ((csa_tree_add_86_2_n_269
    & csa_tree_add_86_2_n_237) | (csa_tree_add_86_2_n_237 & csa_tree_add_86_2_n_327)));
 assign csa_tree_add_86_2_n_545 = (csa_tree_add_86_2_n_269 ^ (csa_tree_add_86_2_n_237 ^ csa_tree_add_86_2_n_327));
 assign csa_tree_add_86_2_n_542 = ((csa_tree_add_86_2_n_356 & csa_tree_add_86_2_n_307) | ((csa_tree_add_86_2_n_307
    & csa_tree_add_86_2_n_244) | (csa_tree_add_86_2_n_244 & csa_tree_add_86_2_n_356)));
 assign csa_tree_add_86_2_n_543 = (csa_tree_add_86_2_n_307 ^ (csa_tree_add_86_2_n_244 ^ csa_tree_add_86_2_n_356));
 assign csa_tree_add_86_2_n_540 = ((csa_tree_add_86_2_n_357 & csa_tree_add_86_2_n_304) | ((csa_tree_add_86_2_n_304
    & csa_tree_add_86_2_n_292) | (csa_tree_add_86_2_n_292 & csa_tree_add_86_2_n_357)));
 assign csa_tree_add_86_2_n_541 = (csa_tree_add_86_2_n_304 ^ (csa_tree_add_86_2_n_292 ^ csa_tree_add_86_2_n_357));
 assign csa_tree_add_86_2_n_538 = ((csa_tree_add_86_2_n_323 & csa_tree_add_86_2_n_305) | ((csa_tree_add_86_2_n_305
    & csa_tree_add_86_2_n_217) | (csa_tree_add_86_2_n_217 & csa_tree_add_86_2_n_323)));
 assign csa_tree_add_86_2_n_539 = (csa_tree_add_86_2_n_305 ^ (csa_tree_add_86_2_n_217 ^ csa_tree_add_86_2_n_323));
 assign csa_tree_add_86_2_n_536 = ((csa_tree_add_86_2_n_330 & csa_tree_add_86_2_n_265) | ((csa_tree_add_86_2_n_265
    & csa_tree_add_86_2_n_239) | (csa_tree_add_86_2_n_239 & csa_tree_add_86_2_n_330)));
 assign csa_tree_add_86_2_n_537 = (csa_tree_add_86_2_n_265 ^ (csa_tree_add_86_2_n_239 ^ csa_tree_add_86_2_n_330));
 assign csa_tree_add_86_2_n_534 = ((csa_tree_add_86_2_n_398 & csa_tree_add_86_2_n_220) | ((csa_tree_add_86_2_n_220
    & csa_tree_add_86_2_n_245) | (csa_tree_add_86_2_n_245 & csa_tree_add_86_2_n_398)));
 assign csa_tree_add_86_2_n_535 = (csa_tree_add_86_2_n_220 ^ (csa_tree_add_86_2_n_245 ^ csa_tree_add_86_2_n_398));
 assign csa_tree_add_86_2_n_532 = ((csa_tree_add_86_2_n_328 & csa_tree_add_86_2_n_246) | ((csa_tree_add_86_2_n_246
    & csa_tree_add_86_2_n_235) | (csa_tree_add_86_2_n_235 & csa_tree_add_86_2_n_328)));
 assign csa_tree_add_86_2_n_533 = (csa_tree_add_86_2_n_246 ^ (csa_tree_add_86_2_n_235 ^ csa_tree_add_86_2_n_328));
 assign csa_tree_add_86_2_n_530 = ((csa_tree_add_86_2_n_335 & csa_tree_add_86_2_n_312) | ((csa_tree_add_86_2_n_312
    & csa_tree_add_86_2_n_286) | (csa_tree_add_86_2_n_286 & csa_tree_add_86_2_n_335)));
 assign csa_tree_add_86_2_n_531 = (csa_tree_add_86_2_n_312 ^ (csa_tree_add_86_2_n_286 ^ csa_tree_add_86_2_n_335));
 assign csa_tree_add_86_2_n_528 = ((csa_tree_add_86_2_n_346 & csa_tree_add_86_2_n_236) | ((csa_tree_add_86_2_n_236
    & csa_tree_add_86_2_n_283) | (csa_tree_add_86_2_n_283 & csa_tree_add_86_2_n_346)));
 assign csa_tree_add_86_2_n_529 = (csa_tree_add_86_2_n_236 ^ (csa_tree_add_86_2_n_283 ^ csa_tree_add_86_2_n_346));
 assign csa_tree_add_86_2_n_526 = ((csa_tree_add_86_2_n_354 & csa_tree_add_86_2_n_255) | ((csa_tree_add_86_2_n_255
    & csa_tree_add_86_2_n_297) | (csa_tree_add_86_2_n_297 & csa_tree_add_86_2_n_354)));
 assign csa_tree_add_86_2_n_527 = (csa_tree_add_86_2_n_255 ^ (csa_tree_add_86_2_n_297 ^ csa_tree_add_86_2_n_354));
 assign csa_tree_add_86_2_n_524 = ((csa_tree_add_86_2_n_397 & csa_tree_add_86_2_n_294) | ((csa_tree_add_86_2_n_294
    & csa_tree_add_86_2_n_268) | (csa_tree_add_86_2_n_268 & csa_tree_add_86_2_n_397)));
 assign csa_tree_add_86_2_n_525 = (csa_tree_add_86_2_n_294 ^ (csa_tree_add_86_2_n_268 ^ csa_tree_add_86_2_n_397));
 assign csa_tree_add_86_2_n_522 = ((csa_tree_add_86_2_n_321 & csa_tree_add_86_2_n_310) | ((csa_tree_add_86_2_n_310
    & csa_tree_add_86_2_n_288) | (csa_tree_add_86_2_n_288 & csa_tree_add_86_2_n_321)));
 assign csa_tree_add_86_2_n_523 = (csa_tree_add_86_2_n_310 ^ (csa_tree_add_86_2_n_288 ^ csa_tree_add_86_2_n_321));
 assign csa_tree_add_86_2_n_520 = ((csa_tree_add_86_2_n_383 & csa_tree_add_86_2_n_316) | ((csa_tree_add_86_2_n_316
    & csa_tree_add_86_2_n_226) | (csa_tree_add_86_2_n_226 & csa_tree_add_86_2_n_383)));
 assign csa_tree_add_86_2_n_521 = (csa_tree_add_86_2_n_316 ^ (csa_tree_add_86_2_n_226 ^ csa_tree_add_86_2_n_383));
 assign csa_tree_add_86_2_n_518 = ((csa_tree_add_86_2_n_412 & csa_tree_add_86_2_n_117) | ((csa_tree_add_86_2_n_117
    & csa_tree_add_86_2_n_181) | (csa_tree_add_86_2_n_181 & csa_tree_add_86_2_n_412)));
 assign csa_tree_add_86_2_n_519 = (csa_tree_add_86_2_n_117 ^ (csa_tree_add_86_2_n_181 ^ csa_tree_add_86_2_n_412));
 assign csa_tree_add_86_2_n_516 = ((csa_tree_add_86_2_n_400 & csa_tree_add_86_2_n_301) | ((csa_tree_add_86_2_n_301
    & csa_tree_add_86_2_n_291) | (csa_tree_add_86_2_n_291 & csa_tree_add_86_2_n_400)));
 assign csa_tree_add_86_2_n_517 = (csa_tree_add_86_2_n_301 ^ (csa_tree_add_86_2_n_291 ^ csa_tree_add_86_2_n_400));
 assign csa_tree_add_86_2_n_514 = ((csa_tree_add_86_2_n_399 & csa_tree_add_86_2_n_264) | ((csa_tree_add_86_2_n_264
    & csa_tree_add_86_2_n_284) | (csa_tree_add_86_2_n_284 & csa_tree_add_86_2_n_399)));
 assign csa_tree_add_86_2_n_515 = (csa_tree_add_86_2_n_264 ^ (csa_tree_add_86_2_n_284 ^ csa_tree_add_86_2_n_399));
 assign csa_tree_add_86_2_n_512 = ((csa_tree_add_86_2_n_360 & csa_tree_add_86_2_n_253) | ((csa_tree_add_86_2_n_253
    & csa_tree_add_86_2_n_254) | (csa_tree_add_86_2_n_254 & csa_tree_add_86_2_n_360)));
 assign csa_tree_add_86_2_n_513 = (csa_tree_add_86_2_n_253 ^ (csa_tree_add_86_2_n_254 ^ csa_tree_add_86_2_n_360));
 assign csa_tree_add_86_2_n_510 = ((csa_tree_add_86_2_n_332 & csa_tree_add_86_2_n_267) | ((csa_tree_add_86_2_n_267
    & csa_tree_add_86_2_n_270) | (csa_tree_add_86_2_n_270 & csa_tree_add_86_2_n_332)));
 assign csa_tree_add_86_2_n_511 = (csa_tree_add_86_2_n_267 ^ (csa_tree_add_86_2_n_270 ^ csa_tree_add_86_2_n_332));
 assign csa_tree_add_86_2_n_508 = ((csa_tree_add_86_2_n_390 & csa_tree_add_86_2_n_90) | ((csa_tree_add_86_2_n_90
    & csa_tree_add_86_2_n_108) | (csa_tree_add_86_2_n_108 & csa_tree_add_86_2_n_390)));
 assign csa_tree_add_86_2_n_509 = (csa_tree_add_86_2_n_90 ^ (csa_tree_add_86_2_n_108 ^ csa_tree_add_86_2_n_390));
 assign csa_tree_add_86_2_n_506 = ((csa_tree_add_86_2_n_396 & csa_tree_add_86_2_n_276) | ((csa_tree_add_86_2_n_276
    & csa_tree_add_86_2_n_258) | (csa_tree_add_86_2_n_258 & csa_tree_add_86_2_n_396)));
 assign csa_tree_add_86_2_n_507 = (csa_tree_add_86_2_n_276 ^ (csa_tree_add_86_2_n_258 ^ csa_tree_add_86_2_n_396));
 assign csa_tree_add_86_2_n_504 = ((csa_tree_add_86_2_n_347 & csa_tree_add_86_2_n_281) | ((csa_tree_add_86_2_n_281
    & csa_tree_add_86_2_n_279) | (csa_tree_add_86_2_n_279 & csa_tree_add_86_2_n_347)));
 assign csa_tree_add_86_2_n_505 = (csa_tree_add_86_2_n_281 ^ (csa_tree_add_86_2_n_279 ^ csa_tree_add_86_2_n_347));
 assign csa_tree_add_86_2_n_502 = ((csa_tree_add_86_2_n_426 & csa_tree_add_86_2_n_130) | ((csa_tree_add_86_2_n_130
    & csa_tree_add_86_2_n_143) | (csa_tree_add_86_2_n_143 & csa_tree_add_86_2_n_426)));
 assign csa_tree_add_86_2_n_503 = (csa_tree_add_86_2_n_130 ^ (csa_tree_add_86_2_n_143 ^ csa_tree_add_86_2_n_426));
 assign csa_tree_add_86_2_n_500 = ((csa_tree_add_86_2_n_336 & csa_tree_add_86_2_n_266) | ((csa_tree_add_86_2_n_266
    & csa_tree_add_86_2_n_314) | (csa_tree_add_86_2_n_314 & csa_tree_add_86_2_n_336)));
 assign csa_tree_add_86_2_n_501 = (csa_tree_add_86_2_n_266 ^ (csa_tree_add_86_2_n_314 ^ csa_tree_add_86_2_n_336));
 assign csa_tree_add_86_2_n_498 = ((csa_tree_add_86_2_n_348 & csa_tree_add_86_2_n_290) | ((csa_tree_add_86_2_n_290
    & csa_tree_add_86_2_n_241) | (csa_tree_add_86_2_n_241 & csa_tree_add_86_2_n_348)));
 assign csa_tree_add_86_2_n_499 = (csa_tree_add_86_2_n_290 ^ (csa_tree_add_86_2_n_241 ^ csa_tree_add_86_2_n_348));
 assign csa_tree_add_86_2_n_496 = ((csa_tree_add_86_2_n_326 & csa_tree_add_86_2_n_251) | ((csa_tree_add_86_2_n_251
    & csa_tree_add_86_2_n_248) | (csa_tree_add_86_2_n_248 & csa_tree_add_86_2_n_326)));
 assign csa_tree_add_86_2_n_497 = (csa_tree_add_86_2_n_251 ^ (csa_tree_add_86_2_n_248 ^ csa_tree_add_86_2_n_326));
 assign csa_tree_add_86_2_n_494 = ((csa_tree_add_86_2_n_343 & csa_tree_add_86_2_n_275) | ((csa_tree_add_86_2_n_275
    & csa_tree_add_86_2_n_285) | (csa_tree_add_86_2_n_285 & csa_tree_add_86_2_n_343)));
 assign csa_tree_add_86_2_n_495 = (csa_tree_add_86_2_n_275 ^ (csa_tree_add_86_2_n_285 ^ csa_tree_add_86_2_n_343));
 assign csa_tree_add_86_2_n_492 = ((csa_tree_add_86_2_n_362 & csa_tree_add_86_2_n_287) | ((csa_tree_add_86_2_n_287
    & csa_tree_add_86_2_n_306) | (csa_tree_add_86_2_n_306 & csa_tree_add_86_2_n_362)));
 assign csa_tree_add_86_2_n_493 = (csa_tree_add_86_2_n_287 ^ (csa_tree_add_86_2_n_306 ^ csa_tree_add_86_2_n_362));
 assign csa_tree_add_86_2_n_490 = ((csa_tree_add_86_2_n_338 & csa_tree_add_86_2_n_308) | ((csa_tree_add_86_2_n_308
    & csa_tree_add_86_2_n_296) | (csa_tree_add_86_2_n_296 & csa_tree_add_86_2_n_338)));
 assign csa_tree_add_86_2_n_491 = (csa_tree_add_86_2_n_308 ^ (csa_tree_add_86_2_n_296 ^ csa_tree_add_86_2_n_338));
 assign csa_tree_add_86_2_n_488 = ((csa_tree_add_86_2_n_337 & csa_tree_add_86_2_n_299) | ((csa_tree_add_86_2_n_299
    & csa_tree_add_86_2_n_260) | (csa_tree_add_86_2_n_260 & csa_tree_add_86_2_n_337)));
 assign csa_tree_add_86_2_n_489 = (csa_tree_add_86_2_n_299 ^ (csa_tree_add_86_2_n_260 ^ csa_tree_add_86_2_n_337));
 assign csa_tree_add_86_2_n_486 = ((csa_tree_add_86_2_n_342 & csa_tree_add_86_2_n_230) | ((csa_tree_add_86_2_n_230
    & csa_tree_add_86_2_n_282) | (csa_tree_add_86_2_n_282 & csa_tree_add_86_2_n_342)));
 assign csa_tree_add_86_2_n_487 = (csa_tree_add_86_2_n_230 ^ (csa_tree_add_86_2_n_282 ^ csa_tree_add_86_2_n_342));
 assign csa_tree_add_86_2_n_484 = ((csa_tree_add_86_2_n_411 & csa_tree_add_86_2_n_116) | ((csa_tree_add_86_2_n_116
    & csa_tree_add_86_2_n_100) | (csa_tree_add_86_2_n_100 & csa_tree_add_86_2_n_411)));
 assign csa_tree_add_86_2_n_485 = (csa_tree_add_86_2_n_116 ^ (csa_tree_add_86_2_n_100 ^ csa_tree_add_86_2_n_411));
 assign csa_tree_add_86_2_n_482 = ((csa_tree_add_86_2_n_402 & csa_tree_add_86_2_n_293) | ((csa_tree_add_86_2_n_293
    & csa_tree_add_86_2_n_317) | (csa_tree_add_86_2_n_317 & csa_tree_add_86_2_n_402)));
 assign csa_tree_add_86_2_n_483 = (csa_tree_add_86_2_n_293 ^ (csa_tree_add_86_2_n_317 ^ csa_tree_add_86_2_n_402));
 assign csa_tree_add_86_2_n_480 = ((csa_tree_add_86_2_n_392 & csa_tree_add_86_2_n_121) | ((csa_tree_add_86_2_n_121
    & csa_tree_add_86_2_n_69) | (csa_tree_add_86_2_n_69 & csa_tree_add_86_2_n_392)));
 assign csa_tree_add_86_2_n_481 = (csa_tree_add_86_2_n_121 ^ (csa_tree_add_86_2_n_69 ^ csa_tree_add_86_2_n_392));
 assign csa_tree_add_86_2_n_478 = ((csa_tree_add_86_2_n_341 & csa_tree_add_86_2_n_274) | ((csa_tree_add_86_2_n_274
    & csa_tree_add_86_2_n_311) | (csa_tree_add_86_2_n_311 & csa_tree_add_86_2_n_341)));
 assign csa_tree_add_86_2_n_479 = (csa_tree_add_86_2_n_274 ^ (csa_tree_add_86_2_n_311 ^ csa_tree_add_86_2_n_341));
 assign csa_tree_add_86_2_n_476 = ((csa_tree_add_86_2_n_351 & csa_tree_add_86_2_n_224) | ((csa_tree_add_86_2_n_224
    & csa_tree_add_86_2_n_240) | (csa_tree_add_86_2_n_240 & csa_tree_add_86_2_n_351)));
 assign csa_tree_add_86_2_n_477 = (csa_tree_add_86_2_n_224 ^ (csa_tree_add_86_2_n_240 ^ csa_tree_add_86_2_n_351));
 assign csa_tree_add_86_2_n_474 = ((csa_tree_add_86_2_n_334 & csa_tree_add_86_2_n_272) | ((csa_tree_add_86_2_n_272
    & csa_tree_add_86_2_n_313) | (csa_tree_add_86_2_n_313 & csa_tree_add_86_2_n_334)));
 assign csa_tree_add_86_2_n_475 = (csa_tree_add_86_2_n_272 ^ (csa_tree_add_86_2_n_313 ^ csa_tree_add_86_2_n_334));
 assign csa_tree_add_86_2_n_472 = ((csa_tree_add_86_2_n_352 & csa_tree_add_86_2_n_300) | ((csa_tree_add_86_2_n_300
    & csa_tree_add_86_2_n_219) | (csa_tree_add_86_2_n_219 & csa_tree_add_86_2_n_352)));
 assign csa_tree_add_86_2_n_473 = (csa_tree_add_86_2_n_300 ^ (csa_tree_add_86_2_n_219 ^ csa_tree_add_86_2_n_352));
 assign csa_tree_add_86_2_n_470 = ((csa_tree_add_86_2_n_202 & csa_tree_add_86_2_n_165) | ((csa_tree_add_86_2_n_165
    & csa_tree_add_86_2_n_152) | (csa_tree_add_86_2_n_152 & csa_tree_add_86_2_n_202)));
 assign csa_tree_add_86_2_n_471 = (csa_tree_add_86_2_n_165 ^ (csa_tree_add_86_2_n_152 ^ csa_tree_add_86_2_n_202));
 assign csa_tree_add_86_2_n_468 = ((csa_tree_add_86_2_n_325 & csa_tree_add_86_2_n_318) | ((csa_tree_add_86_2_n_318
    & csa_tree_add_86_2_n_309) | (csa_tree_add_86_2_n_309 & csa_tree_add_86_2_n_325)));
 assign csa_tree_add_86_2_n_469 = (csa_tree_add_86_2_n_318 ^ (csa_tree_add_86_2_n_309 ^ csa_tree_add_86_2_n_325));
 assign csa_tree_add_86_2_n_466 = ((csa_tree_add_86_2_n_333 & csa_tree_add_86_2_n_315) | ((csa_tree_add_86_2_n_315
    & csa_tree_add_86_2_n_280) | (csa_tree_add_86_2_n_280 & csa_tree_add_86_2_n_333)));
 assign csa_tree_add_86_2_n_467 = (csa_tree_add_86_2_n_315 ^ (csa_tree_add_86_2_n_280 ^ csa_tree_add_86_2_n_333));
 assign csa_tree_add_86_2_n_462 = ((csa_tree_add_86_2_n_212 & csa_tree_add_86_2_n_104) | ((csa_tree_add_86_2_n_104
    & csa_tree_add_86_2_n_38) | (csa_tree_add_86_2_n_38 & csa_tree_add_86_2_n_212)));
 assign csa_tree_add_86_2_n_463 = (csa_tree_add_86_2_n_104 ^ (csa_tree_add_86_2_n_38 ^ csa_tree_add_86_2_n_212));
 assign csa_tree_add_86_2_n_460 = ((csa_tree_add_86_2_n_339 & csa_tree_add_86_2_n_242) | ((csa_tree_add_86_2_n_242
    & csa_tree_add_86_2_n_225) | (csa_tree_add_86_2_n_225 & csa_tree_add_86_2_n_339)));
 assign csa_tree_add_86_2_n_461 = (csa_tree_add_86_2_n_242 ^ (csa_tree_add_86_2_n_225 ^ csa_tree_add_86_2_n_339));
 assign csa_tree_add_86_2_n_458 = ((csa_tree_add_86_2_n_324 & csa_tree_add_86_2_n_273) | ((csa_tree_add_86_2_n_273
    & csa_tree_add_86_2_n_234) | (csa_tree_add_86_2_n_234 & csa_tree_add_86_2_n_324)));
 assign csa_tree_add_86_2_n_459 = (csa_tree_add_86_2_n_273 ^ (csa_tree_add_86_2_n_234 ^ csa_tree_add_86_2_n_324));
 assign csa_tree_add_86_2_n_456 = ((csa_tree_add_86_2_n_194 & csa_tree_add_86_2_n_146) | ((csa_tree_add_86_2_n_146
    & csa_tree_add_86_2_n_221) | (csa_tree_add_86_2_n_221 & csa_tree_add_86_2_n_194)));
 assign csa_tree_add_86_2_n_457 = (csa_tree_add_86_2_n_146 ^ (csa_tree_add_86_2_n_221 ^ csa_tree_add_86_2_n_194));
 assign csa_tree_add_86_2_n_454 = ((csa_tree_add_86_2_n_208 & csa_tree_add_86_2_n_183) | ((csa_tree_add_86_2_n_183
    & csa_tree_add_86_2_n_113) | (csa_tree_add_86_2_n_113 & csa_tree_add_86_2_n_208)));
 assign csa_tree_add_86_2_n_455 = (csa_tree_add_86_2_n_183 ^ (csa_tree_add_86_2_n_113 ^ csa_tree_add_86_2_n_208));
 assign csa_tree_add_86_2_n_452 = ((csa_tree_add_86_2_n_320 & csa_tree_add_86_2_n_177) | ((csa_tree_add_86_2_n_177
    & csa_tree_add_86_2_n_118) | (csa_tree_add_86_2_n_118 & csa_tree_add_86_2_n_320)));
 assign csa_tree_add_86_2_n_453 = (csa_tree_add_86_2_n_177 ^ (csa_tree_add_86_2_n_118 ^ csa_tree_add_86_2_n_320));
 assign csa_tree_add_86_2_n_450 = ((csa_tree_add_86_2_n_204 & csa_tree_add_86_2_n_167) | ((csa_tree_add_86_2_n_167
    & csa_tree_add_86_2_n_51) | (csa_tree_add_86_2_n_51 & csa_tree_add_86_2_n_204)));
 assign csa_tree_add_86_2_n_451 = (csa_tree_add_86_2_n_167 ^ (csa_tree_add_86_2_n_51 ^ csa_tree_add_86_2_n_204));
 assign csa_tree_add_86_2_n_448 = ((csa_tree_add_86_2_n_363 & csa_tree_add_86_2_n_87) | ((csa_tree_add_86_2_n_87
    & csa_tree_add_86_2_n_142) | (csa_tree_add_86_2_n_142 & csa_tree_add_86_2_n_363)));
 assign csa_tree_add_86_2_n_449 = (csa_tree_add_86_2_n_87 ^ (csa_tree_add_86_2_n_142 ^ csa_tree_add_86_2_n_363));
 assign csa_tree_add_86_2_n_446 = ((csa_tree_add_86_2_n_210 & csa_tree_add_86_2_n_99) | ((csa_tree_add_86_2_n_99
    & csa_tree_add_86_2_n_65) | (csa_tree_add_86_2_n_65 & csa_tree_add_86_2_n_210)));
 assign csa_tree_add_86_2_n_447 = (csa_tree_add_86_2_n_99 ^ (csa_tree_add_86_2_n_65 ^ csa_tree_add_86_2_n_210));
 assign csa_tree_add_86_2_n_444 = ((csa_tree_add_86_2_n_196 & csa_tree_add_86_2_n_252) | ((csa_tree_add_86_2_n_252
    & csa_tree_add_86_2_n_289) | (csa_tree_add_86_2_n_289 & csa_tree_add_86_2_n_196)));
 assign csa_tree_add_86_2_n_445 = (csa_tree_add_86_2_n_252 ^ (csa_tree_add_86_2_n_289 ^ csa_tree_add_86_2_n_196));
 assign csa_tree_add_86_2_n_442 = ((csa_tree_add_86_2_n_197 & csa_tree_add_86_2_n_271) | ((csa_tree_add_86_2_n_271
    & csa_tree_add_86_2_n_302) | (csa_tree_add_86_2_n_302 & csa_tree_add_86_2_n_197)));
 assign csa_tree_add_86_2_n_443 = (csa_tree_add_86_2_n_271 ^ (csa_tree_add_86_2_n_302 ^ csa_tree_add_86_2_n_197));
 assign csa_tree_add_86_2_n_440 = ((csa_tree_add_86_2_n_195 & csa_tree_add_86_2_n_190) | ((csa_tree_add_86_2_n_190
    & csa_tree_add_86_2_n_247) | (csa_tree_add_86_2_n_247 & csa_tree_add_86_2_n_195)));
 assign csa_tree_add_86_2_n_441 = (csa_tree_add_86_2_n_190 ^ (csa_tree_add_86_2_n_247 ^ csa_tree_add_86_2_n_195));
 assign csa_tree_add_86_2_n_438 = ((csa_tree_add_86_2_n_211 & csa_tree_add_86_2_n_55) | ((csa_tree_add_86_2_n_55
    & csa_tree_add_86_2_n_119) | (csa_tree_add_86_2_n_119 & csa_tree_add_86_2_n_211)));
 assign csa_tree_add_86_2_n_439 = (csa_tree_add_86_2_n_55 ^ (csa_tree_add_86_2_n_119 ^ csa_tree_add_86_2_n_211));
 assign csa_tree_add_86_2_n_436 = ((csa_tree_add_86_2_n_207 & csa_tree_add_86_2_n_58) | ((csa_tree_add_86_2_n_58
    & csa_tree_add_86_2_n_148) | (csa_tree_add_86_2_n_148 & csa_tree_add_86_2_n_207)));
 assign csa_tree_add_86_2_n_437 = (csa_tree_add_86_2_n_58 ^ (csa_tree_add_86_2_n_148 ^ csa_tree_add_86_2_n_207));
 assign csa_tree_add_86_2_n_434 = ((csa_tree_add_86_2_n_377 & csa_tree_add_86_2_n_159) | ((csa_tree_add_86_2_n_159
    & csa_tree_add_86_2_n_178) | (csa_tree_add_86_2_n_178 & csa_tree_add_86_2_n_377)));
 assign csa_tree_add_86_2_n_435 = (csa_tree_add_86_2_n_159 ^ (csa_tree_add_86_2_n_178 ^ csa_tree_add_86_2_n_377));
 assign csa_tree_add_86_2_n_430 = ((csa_tree_add_86_2_n_322 & csa_tree_add_86_2_n_259) | ((csa_tree_add_86_2_n_259
    & csa_tree_add_86_2_n_228) | (csa_tree_add_86_2_n_228 & csa_tree_add_86_2_n_322)));
 assign csa_tree_add_86_2_n_431 = (csa_tree_add_86_2_n_259 ^ (csa_tree_add_86_2_n_228 ^ csa_tree_add_86_2_n_322));
 assign csa_tree_add_86_2_n_428 = ((csa_tree_add_86_2_n_384 & csa_tree_add_86_2_n_145) | ((csa_tree_add_86_2_n_145
    & csa_tree_add_86_2_n_114) | (csa_tree_add_86_2_n_114 & csa_tree_add_86_2_n_384)));
 assign csa_tree_add_86_2_n_429 = (csa_tree_add_86_2_n_145 ^ (csa_tree_add_86_2_n_114 ^ csa_tree_add_86_2_n_384));
 assign csa_tree_add_86_2_n_426 = (csa_tree_add_86_2_n_199 & csa_tree_add_86_2_n_373);
 assign csa_tree_add_86_2_n_427 = (csa_tree_add_86_2_n_199 ^ csa_tree_add_86_2_n_373);
 assign csa_tree_add_86_2_n_424 = (csa_tree_add_86_2_n_372 & csa_tree_add_86_2_n_374);
 assign csa_tree_add_86_2_n_425 = (csa_tree_add_86_2_n_372 ^ csa_tree_add_86_2_n_374);
 assign csa_tree_add_86_2_n_422 = (csa_tree_add_86_2_n_193 & csa_tree_add_86_2_n_366);
 assign csa_tree_add_86_2_n_423 = (csa_tree_add_86_2_n_193 ^ csa_tree_add_86_2_n_366);
 assign csa_tree_add_86_2_n_420 = (csa_tree_add_86_2_n_369 & csa_tree_add_86_2_n_355);
 assign csa_tree_add_86_2_n_421 = (csa_tree_add_86_2_n_369 ^ csa_tree_add_86_2_n_355);
 assign csa_tree_add_86_2_n_418 = (csa_tree_add_86_2_n_319 & csa_tree_add_86_2_n_365);
 assign csa_tree_add_86_2_n_419 = (csa_tree_add_86_2_n_319 ^ csa_tree_add_86_2_n_365);
 assign csa_tree_add_86_2_n_416 = (csa_tree_add_86_2_n_203 & csa_tree_add_86_2_n_381);
 assign csa_tree_add_86_2_n_417 = (csa_tree_add_86_2_n_203 ^ csa_tree_add_86_2_n_381);
 assign csa_tree_add_86_2_n_414 = (csa_tree_add_86_2_n_205 & csa_tree_add_86_2_n_379);
 assign csa_tree_add_86_2_n_415 = (csa_tree_add_86_2_n_205 ^ csa_tree_add_86_2_n_379);
 assign csa_tree_add_86_2_n_412 = (csa_tree_add_86_2_n_200 & csa_tree_add_86_2_n_368);
 assign csa_tree_add_86_2_n_413 = (csa_tree_add_86_2_n_200 ^ csa_tree_add_86_2_n_368);
 assign csa_tree_add_86_2_n_410 = (csa_tree_add_86_2_n_385 & csa_tree_add_86_2_n_361);
 assign csa_tree_add_86_2_n_411 = (csa_tree_add_86_2_n_385 ^ csa_tree_add_86_2_n_361);
 assign csa_tree_add_86_2_n_408 = (csa_tree_add_86_2_n_206 & csa_tree_add_86_2_n_378);
 assign csa_tree_add_86_2_n_409 = (csa_tree_add_86_2_n_206 ^ csa_tree_add_86_2_n_378);
 assign csa_tree_add_86_2_n_406 = (csa_tree_add_86_2_n_387 & csa_tree_add_86_2_n_370);
 assign csa_tree_add_86_2_n_407 = (csa_tree_add_86_2_n_387 ^ csa_tree_add_86_2_n_370);
 assign csa_tree_add_86_2_n_404 = (csa_tree_add_86_2_n_344 & csa_tree_add_86_2_n_353);
 assign csa_tree_add_86_2_n_405 = (csa_tree_add_86_2_n_344 ^ csa_tree_add_86_2_n_353);
 assign csa_tree_add_86_2_n_402 = (csa_tree_add_86_2_n_349 & csa_tree_add_86_2_n_340);
 assign csa_tree_add_86_2_n_403 = (csa_tree_add_86_2_n_349 ^ csa_tree_add_86_2_n_340);
 assign csa_tree_add_86_2_n_400 = (csa_tree_add_86_2_n_371 & csa_tree_add_86_2_n_358);
 assign n_1377 = (csa_tree_add_86_2_n_371 ^ csa_tree_add_86_2_n_358);
 assign csa_tree_add_86_2_n_398 = (csa_tree_add_86_2_n_329 & csa_tree_add_86_2_n_331);
 assign csa_tree_add_86_2_n_399 = (csa_tree_add_86_2_n_329 ^ csa_tree_add_86_2_n_331);
 assign csa_tree_add_86_2_n_396 = (csa_tree_add_86_2_n_359 & csa_tree_add_86_2_n_364);
 assign csa_tree_add_86_2_n_397 = (csa_tree_add_86_2_n_359 ^ csa_tree_add_86_2_n_364);
 assign csa_tree_add_86_2_n_394 = (csa_tree_add_86_2_n_201 & csa_tree_add_86_2_n_375);
 assign csa_tree_add_86_2_n_395 = (csa_tree_add_86_2_n_201 ^ csa_tree_add_86_2_n_375);
 assign csa_tree_add_86_2_n_392 = (csa_tree_add_86_2_n_209 & csa_tree_add_86_2_n_376);
 assign csa_tree_add_86_2_n_393 = (csa_tree_add_86_2_n_209 ^ csa_tree_add_86_2_n_376);
 assign csa_tree_add_86_2_n_390 = (csa_tree_add_86_2_n_213 & csa_tree_add_86_2_n_367);
 assign csa_tree_add_86_2_n_391 = (csa_tree_add_86_2_n_213 ^ csa_tree_add_86_2_n_367);
 assign csa_tree_add_86_2_n_388 = (csa_tree_add_86_2_n_386 & csa_tree_add_86_2_n_380);
 assign csa_tree_add_86_2_n_389 = (csa_tree_add_86_2_n_386 ^ csa_tree_add_86_2_n_380);
 assign csa_tree_add_86_2_n_383 = ({in3[6]} & {in4[6]});
 assign csa_tree_add_86_2_n_382 = ~(csa_tree_add_86_2_n_28 | csa_tree_add_86_2_n_31);
 assign csa_tree_add_86_2_n_374 = ({in1[0]} & {in2[4]});
 assign csa_tree_add_86_2_n_372 = ({in3[4]} & {in4[0]});
 assign csa_tree_add_86_2_n_371 = ({in3[0]} & {in4[0]});
 assign csa_tree_add_86_2_n_369 = ({in3[6]} & {in4[0]});
 assign csa_tree_add_86_2_n_365 = ({in1[1]} & {in2[4]});
 assign csa_tree_add_86_2_n_364 = ({in1[4]} & {in2[6]});
 assign csa_tree_add_86_2_n_362 = ({in3[7]} & {in4[5]});
 assign csa_tree_add_86_2_n_360 = ({in3[3]} & {in4[6]});
 assign csa_tree_add_86_2_n_359 = ({in1[3]} & {in2[7]});
 assign csa_tree_add_86_2_n_358 = ({in1[0]} & {in2[0]});
 assign csa_tree_add_86_2_n_357 = ({in1[4]} & {in2[5]});
 assign csa_tree_add_86_2_n_356 = ({in3[3]} & {in4[3]});
 assign csa_tree_add_86_2_n_355 = ({in1[0]} & {in2[6]});
 assign csa_tree_add_86_2_n_354 = ({in3[0]} & {in4[5]});
 assign csa_tree_add_86_2_n_353 = ({in1[1]} & {in2[0]});
 assign csa_tree_add_86_2_n_352 = ({in1[5]} & {in2[3]});
 assign csa_tree_add_86_2_n_351 = ({in1[6]} & {in2[5]});
 assign csa_tree_add_86_2_n_350 = ({in3[1]} & {in4[1]});
 assign csa_tree_add_86_2_n_349 = ({in1[0]} & {in2[3]});
 assign csa_tree_add_86_2_n_348 = ({in1[4]} & {in2[2]});
 assign csa_tree_add_86_2_n_347 = ({in3[6]} & {in4[4]});
 assign csa_tree_add_86_2_n_346 = ({in3[4]} & {in4[3]});
 assign csa_tree_add_86_2_n_345 = ({in3[2]} & {in4[2]});
 assign csa_tree_add_86_2_n_344 = ({in1[0]} & {in2[1]});
 assign csa_tree_add_86_2_n_343 = ({in1[2]} & {in2[5]});
 assign csa_tree_add_86_2_n_342 = ({in3[5]} & {in4[0]});
 assign csa_tree_add_86_2_n_341 = ({in1[1]} & {in2[1]});
 assign csa_tree_add_86_2_n_340 = ({in1[3]} & {in2[0]});
 assign csa_tree_add_86_2_n_338 = ({in3[1]} & {in4[2]});
 assign csa_tree_add_86_2_n_337 = ({in1[6]} & {in2[0]});
 assign csa_tree_add_86_2_n_336 = ({in3[7]} & {in4[3]});
 assign csa_tree_add_86_2_n_335 = ({in1[5]} & {in2[4]});
 assign csa_tree_add_86_2_n_334 = ({in1[5]} & {in2[6]});
 assign csa_tree_add_86_2_n_333 = ({in1[7]} & {in2[6]});
 assign csa_tree_add_86_2_n_332 = ({in3[4]} & {in4[1]});
 assign csa_tree_add_86_2_n_331 = ({in1[1]} & {in2[6]});
 assign csa_tree_add_86_2_n_330 = ({in3[7]} & {in4[2]});
 assign csa_tree_add_86_2_n_329 = ({in1[0]} & {in2[7]});
 assign csa_tree_add_86_2_n_328 = ({in3[1]} & {in4[6]});
 assign csa_tree_add_86_2_n_327 = ({in1[2]} & {in2[1]});
 assign csa_tree_add_86_2_n_326 = ({in1[4]} & {in2[0]});
 assign csa_tree_add_86_2_n_325 = ({in3[6]} & {in4[2]});
 assign csa_tree_add_86_2_n_324 = ({in3[3]} & {in4[5]});
 assign csa_tree_add_86_2_n_323 = ({in3[6]} & {in4[1]});
 assign csa_tree_add_86_2_n_322 = ({in1[2]} & {in2[6]});
 assign csa_tree_add_86_2_n_321 = ({in1[1]} & {in2[5]});
 assign csa_tree_add_86_2_n_319 = ({in1[0]} & {in2[5]});
 assign csa_tree_add_86_2_n_318 = ({in1[7]} & {in2[1]});
 assign csa_tree_add_86_2_n_317 = ({in3[3]} & {in4[1]});
 assign csa_tree_add_86_2_n_316 = ({in1[6]} & {in2[6]});
 assign csa_tree_add_86_2_n_315 = ({in3[6]} & {in4[7]});
 assign csa_tree_add_86_2_n_314 = ({in3[5]} & {in4[5]});
 assign csa_tree_add_86_2_n_313 = ({in3[5]} & {in4[6]});
 assign csa_tree_add_86_2_n_312 = ({in3[4]} & {in4[5]});
 assign csa_tree_add_86_2_n_311 = ({in3[0]} & {in4[2]});
 assign csa_tree_add_86_2_n_310 = ({in3[4]} & {in4[2]});
 assign csa_tree_add_86_2_n_309 = ({in3[7]} & {in4[1]});
 assign csa_tree_add_86_2_n_308 = ({in1[1]} & {in2[2]});
 assign csa_tree_add_86_2_n_307 = ({in3[5]} & {in4[1]});
 assign csa_tree_add_86_2_n_306 = ({in3[5]} & {in4[7]});
 assign csa_tree_add_86_2_n_305 = ({in1[6]} & {in2[1]});
 assign csa_tree_add_86_2_n_304 = ({in1[3]} & {in2[6]});
 assign csa_tree_add_86_2_n_303 = ({in1[5]} & {in2[0]});
 assign csa_tree_add_86_2_n_301 = ({in3[1]} & {in4[0]});
 assign csa_tree_add_86_2_n_300 = ({in1[6]} & {in2[2]});
 assign csa_tree_add_86_2_n_299 = ({in1[3]} & {in2[3]});
 assign csa_tree_add_86_2_n_297 = ({in3[1]} & {in4[4]});
 assign csa_tree_add_86_2_n_296 = ({in3[3]} & {in4[0]});
 assign csa_tree_add_86_2_n_294 = ({in3[4]} & {in4[6]});
 assign csa_tree_add_86_2_n_293 = ({in1[3]} & {in2[1]});
 assign csa_tree_add_86_2_n_292 = ({in1[2]} & {in2[7]});
 assign csa_tree_add_86_2_n_291 = ({in3[0]} & {in4[1]});
 assign csa_tree_add_86_2_n_290 = ({in1[5]} & {in2[1]});
 assign csa_tree_add_86_2_n_288 = ({in3[1]} & {in4[5]});
 assign csa_tree_add_86_2_n_287 = ({in1[7]} & {in2[5]});
 assign csa_tree_add_86_2_n_286 = ({in3[2]} & {in4[7]});
 assign csa_tree_add_86_2_n_285 = ({in3[7]} & {in4[0]});
 assign csa_tree_add_86_2_n_284 = ({in3[0]} & {in4[7]});
 assign csa_tree_add_86_2_n_283 = ({in1[3]} & {in2[4]});
 assign csa_tree_add_86_2_n_282 = ({in3[2]} & {in4[3]});
 assign csa_tree_add_86_2_n_281 = ({in1[7]} & {in2[3]});
 assign csa_tree_add_86_2_n_280 = ({in1[6]} & {in2[7]});
 assign csa_tree_add_86_2_n_279 = ({in1[5]} & {in2[5]});
 assign csa_tree_add_86_2_n_278 = ({in3[1]} & {in4[3]});
 assign csa_tree_add_86_2_n_276 = ({in1[7]} & {in2[4]});
 assign csa_tree_add_86_2_n_275 = ({in1[7]} & {in2[0]});
 assign csa_tree_add_86_2_n_274 = ({in1[2]} & {in2[0]});
 assign csa_tree_add_86_2_n_273 = ({in1[4]} & {in2[4]});
 assign csa_tree_add_86_2_n_272 = ({in1[4]} & {in2[7]});
 assign csa_tree_add_86_2_n_270 = ({in1[2]} & {in2[3]});
 assign csa_tree_add_86_2_n_269 = ({in3[2]} & {in4[1]});
 assign csa_tree_add_86_2_n_268 = ({in3[3]} & {in4[7]});
 assign csa_tree_add_86_2_n_267 = ({in1[4]} & {in2[1]});
 assign csa_tree_add_86_2_n_266 = ({in1[6]} & {in2[4]});
 assign csa_tree_add_86_2_n_265 = ({in1[6]} & {in2[3]});
 assign csa_tree_add_86_2_n_264 = ({in3[5]} & {in4[2]});
 assign csa_tree_add_86_2_n_263 = ({in3[7]} & {in4[6]});
 assign csa_tree_add_86_2_n_262 = ({in3[2]} & {in4[0]});
 assign csa_tree_add_86_2_n_261 = ({in1[0]} & {in2[2]});
 assign csa_tree_add_86_2_n_260 = ({in3[0]} & {in4[6]});
 assign csa_tree_add_86_2_n_259 = ({in1[3]} & {in2[5]});
 assign csa_tree_add_86_2_n_258 = ({in3[6]} & {in4[5]});
 assign csa_tree_add_86_2_n_257 = ({in3[0]} & {in4[4]});
 assign csa_tree_add_86_2_n_256 = ({in3[7]} & {in4[7]});
 assign csa_tree_add_86_2_n_255 = ({in1[3]} & {in2[2]});
 assign csa_tree_add_86_2_n_254 = ({in3[5]} & {in4[4]});
 assign csa_tree_add_86_2_n_253 = ({in1[7]} & {in2[2]});
 assign csa_tree_add_86_2_n_251 = ({in1[2]} & {in2[2]});
 assign csa_tree_add_86_2_n_250 = ~(csa_tree_add_86_2_n_29 | csa_tree_add_86_2_n_21);
 assign csa_tree_add_86_2_n_249 = ~(csa_tree_add_86_2_n_29 | csa_tree_add_86_2_n_11);
 assign csa_tree_add_86_2_n_248 = ({in1[1]} & {in2[3]});
 assign csa_tree_add_86_2_n_246 = ({in3[3]} & {in4[4]});
 assign csa_tree_add_86_2_n_245 = ({in3[4]} & {in4[4]});
 assign csa_tree_add_86_2_n_244 = ({in3[2]} & {in4[4]});
 assign csa_tree_add_86_2_n_243 = ~(csa_tree_add_86_2_n_29 | csa_tree_add_86_2_n_31);
 assign csa_tree_add_86_2_n_241 = ({in1[2]} & {in2[4]});
 assign csa_tree_add_86_2_n_240 = ({in3[7]} & {in4[4]});
 assign csa_tree_add_86_2_n_239 = ({in3[6]} & {in4[3]});
 assign csa_tree_add_86_2_n_238 = ~(csa_tree_add_86_2_n_29 | csa_tree_add_86_2_n_33);
 assign csa_tree_add_86_2_n_237 = ({in3[0]} & {in4[3]});
 assign csa_tree_add_86_2_n_236 = ({in1[4]} & {in2[3]});
 assign csa_tree_add_86_2_n_235 = ({in3[2]} & {in4[5]});
 assign csa_tree_add_86_2_n_234 = ({in3[2]} & {in4[6]});
 assign csa_tree_add_86_2_n_233 = ~(csa_tree_add_86_2_n_29 | csa_tree_add_86_2_n_12);
 assign csa_tree_add_86_2_n_232 = ~(csa_tree_add_86_2_n_29 | csa_tree_add_86_2_n_18);
 assign csa_tree_add_86_2_n_231 = ~(csa_tree_add_86_2_n_29 | csa_tree_add_86_2_n_20);
 assign csa_tree_add_86_2_n_230 = ({in3[3]} & {in4[2]});
 assign csa_tree_add_86_2_n_229 = ~(csa_tree_add_86_2_n_29 | csa_tree_add_86_2_n_35);
 assign csa_tree_add_86_2_n_228 = ({in1[1]} & {in2[7]});
 assign csa_tree_add_86_2_n_227 = ~(csa_tree_add_86_2_n_29 | csa_tree_add_86_2_n_37);
 assign csa_tree_add_86_2_n_226 = ({in1[5]} & {in2[7]});
 assign csa_tree_add_86_2_n_224 = ({in3[4]} & {in4[7]});
 assign csa_tree_add_86_2_n_223 = ~(csa_tree_add_86_2_n_28 | csa_tree_add_86_2_n_11);
 assign csa_tree_add_86_2_n_222 = ~(csa_tree_add_86_2_n_28 | csa_tree_add_86_2_n_21);
 assign csa_tree_add_86_2_n_220 = ({in3[5]} & {in4[3]});
 assign csa_tree_add_86_2_n_219 = ({in3[1]} & {in4[7]});
 assign csa_tree_add_86_2_n_218 = ({in1[7]} & {in2[7]});
 assign csa_tree_add_86_2_n_217 = ({in1[5]} & {in2[2]});
 assign n_1407 = ~(csa_tree_add_86_2_n_5 | csa_tree_add_86_2_n_11);
 assign n_1376 = ~(csa_tree_add_86_2_n_5 | csa_tree_add_86_2_n_37);
 assign n_1375 = ~(csa_tree_add_86_2_n_5 | csa_tree_add_86_2_n_20);
 assign csa_tree_add_86_2_n_207 = ~(csa_tree_add_86_2_n_4 | csa_tree_add_86_2_n_18);
 assign csa_tree_add_86_2_n_198 = ~(csa_tree_add_86_2_n_27 | csa_tree_add_86_2_n_18);
 assign csa_tree_add_86_2_n_192 = ~(csa_tree_add_86_2_n_3 | csa_tree_add_86_2_n_18);
 assign csa_tree_add_86_2_n_189 = ~(csa_tree_add_86_2_n_3 | csa_tree_add_86_2_n_11);
 assign csa_tree_add_86_2_n_188 = ~(csa_tree_add_86_2_n_3 | csa_tree_add_86_2_n_12);
 assign csa_tree_add_86_2_n_186 = ({in5[0]} & n_1341);
 assign csa_tree_add_86_2_n_184 = ~(csa_tree_add_86_2_n_26 | csa_tree_add_86_2_n_37);
 assign csa_tree_add_86_2_n_182 = ~(csa_tree_add_86_2_n_28 | csa_tree_add_86_2_n_12);
 assign csa_tree_add_86_2_n_179 = ~(csa_tree_add_86_2_n_5 | csa_tree_add_86_2_n_35);
 assign csa_tree_add_86_2_n_175 = ~(csa_tree_add_86_2_n_3 | csa_tree_add_86_2_n_33);
 assign csa_tree_add_86_2_n_174 = ~(csa_tree_add_86_2_n_27 | csa_tree_add_86_2_n_12);
 assign csa_tree_add_86_2_n_173 = ~(csa_tree_add_86_2_n_4 | csa_tree_add_86_2_n_31);
 assign csa_tree_add_86_2_n_172 = ~(csa_tree_add_86_2_n_5 | csa_tree_add_86_2_n_33);
 assign csa_tree_add_86_2_n_171 = ~(csa_tree_add_86_2_n_4 | csa_tree_add_86_2_n_11);
 assign csa_tree_add_86_2_n_169 = ~(csa_tree_add_86_2_n_28 | csa_tree_add_86_2_n_33);
 assign csa_tree_add_86_2_n_166 = ({in5[1]} & n_1496);
 assign csa_tree_add_86_2_n_164 = ~(csa_tree_add_86_2_n_25 | csa_tree_add_86_2_n_31);
 assign csa_tree_add_86_2_n_162 = ~(csa_tree_add_86_2_n_27 | csa_tree_add_86_2_n_33);
 assign csa_tree_add_86_2_n_161 = ~(csa_tree_add_86_2_n_28 | csa_tree_add_86_2_n_20);
 assign csa_tree_add_86_2_n_158 = ({in5[0]} & n_1339);
 assign csa_tree_add_86_2_n_157 = ~(csa_tree_add_86_2_n_4 | csa_tree_add_86_2_n_33);
 assign csa_tree_add_86_2_n_156 = ~(csa_tree_add_86_2_n_26 | csa_tree_add_86_2_n_6);
 assign csa_tree_add_86_2_n_154 = ~(csa_tree_add_86_2_n_28 | csa_tree_add_86_2_n_18);
 assign csa_tree_add_86_2_n_153 = ~(csa_tree_add_86_2_n_25 | csa_tree_add_86_2_n_37);
 assign csa_tree_add_86_2_n_151 = ~(csa_tree_add_86_2_n_25 | csa_tree_add_86_2_n_18);
 assign csa_tree_add_86_2_n_148 = ~(csa_tree_add_86_2_n_25 | n_1498);
 assign csa_tree_add_86_2_n_147 = ~(csa_tree_add_86_2_n_25 | csa_tree_add_86_2_n_35);
 assign csa_tree_add_86_2_n_144 = ~(csa_tree_add_86_2_n_26 | csa_tree_add_86_2_n_20);
 assign csa_tree_add_86_2_n_141 = ~(csa_tree_add_86_2_n_26 | n_1498);
 assign csa_tree_add_86_2_n_140 = ~(csa_tree_add_86_2_n_27 | csa_tree_add_86_2_n_20);
 assign csa_tree_add_86_2_n_139 = ({in5[0]} & n_1340);
 assign csa_tree_add_86_2_n_133 = ~(csa_tree_add_86_2_n_26 | csa_tree_add_86_2_n_35);
 assign csa_tree_add_86_2_n_132 = ~(csa_tree_add_86_2_n_25 | csa_tree_add_86_2_n_7);
 assign csa_tree_add_86_2_n_131 = ~(csa_tree_add_86_2_n_5 | csa_tree_add_86_2_n_21);
 assign csa_tree_add_86_2_n_127 = ~(csa_tree_add_86_2_n_28 | csa_tree_add_86_2_n_35);
 assign csa_tree_add_86_2_n_126 = ~(csa_tree_add_86_2_n_28 | csa_tree_add_86_2_n_37);
 assign csa_tree_add_86_2_n_125 = ~(csa_tree_add_86_2_n_4 | n_1498);
 assign csa_tree_add_86_2_n_122 = ~(csa_tree_add_86_2_n_27 | csa_tree_add_86_2_n_35);
 assign csa_tree_add_86_2_n_111 = ~(csa_tree_add_86_2_n_27 | csa_tree_add_86_2_n_21);
 assign csa_tree_add_86_2_n_109 = ~(csa_tree_add_86_2_n_3 | n_1498);
 assign csa_tree_add_86_2_n_106 = ~(csa_tree_add_86_2_n_25 | csa_tree_add_86_2_n_21);
 assign csa_tree_add_86_2_n_105 = ~(csa_tree_add_86_2_n_27 | n_1498);
 assign csa_tree_add_86_2_n_101 = ~(csa_tree_add_86_2_n_26 | csa_tree_add_86_2_n_21);
 assign csa_tree_add_86_2_n_98 = ~(csa_tree_add_86_2_n_5 | csa_tree_add_86_2_n_18);
 assign csa_tree_add_86_2_n_95 = ~(csa_tree_add_86_2_n_4 | csa_tree_add_86_2_n_37);
 assign csa_tree_add_86_2_n_94 = ~(csa_tree_add_86_2_n_27 | csa_tree_add_86_2_n_37);
 assign csa_tree_add_86_2_n_91 = ~(csa_tree_add_86_2_n_27 | csa_tree_add_86_2_n_11);
 assign csa_tree_add_86_2_n_86 = ~(csa_tree_add_86_2_n_25 | csa_tree_add_86_2_n_33);
 assign csa_tree_add_86_2_n_84 = ~(csa_tree_add_86_2_n_25 | csa_tree_add_86_2_n_11);
 assign csa_tree_add_86_2_n_83 = ~(n_1498 | ~{in5[0]});
 assign csa_tree_add_86_2_n_82 = ~(csa_tree_add_86_2_n_3 | csa_tree_add_86_2_n_37);
 assign csa_tree_add_86_2_n_81 = ~(csa_tree_add_86_2_n_3 | csa_tree_add_86_2_n_31);
 assign csa_tree_add_86_2_n_76 = ({in5[1]} & n_1344);
 assign csa_tree_add_86_2_n_75 = ~(csa_tree_add_86_2_n_25 | csa_tree_add_86_2_n_20);
 assign csa_tree_add_86_2_n_74 = ~(csa_tree_add_86_2_n_4 | csa_tree_add_86_2_n_12);
 assign csa_tree_add_86_2_n_72 = ~(csa_tree_add_86_2_n_26 | csa_tree_add_86_2_n_11);
 assign csa_tree_add_86_2_n_68 = ~(csa_tree_add_86_2_n_3 | csa_tree_add_86_2_n_35);
 assign csa_tree_add_86_2_n_67 = ~(csa_tree_add_86_2_n_5 | csa_tree_add_86_2_n_31);
 assign csa_tree_add_86_2_n_66 = ~(csa_tree_add_86_2_n_5 | csa_tree_add_86_2_n_12);
 assign csa_tree_add_86_2_n_61 = ~(csa_tree_add_86_2_n_26 | csa_tree_add_86_2_n_33);
 assign csa_tree_add_86_2_n_59 = ~(csa_tree_add_86_2_n_4 | csa_tree_add_86_2_n_20);
 assign csa_tree_add_86_2_n_58 = ~(csa_tree_add_86_2_n_26 | csa_tree_add_86_2_n_7);
 assign csa_tree_add_86_2_n_57 = ~(csa_tree_add_86_2_n_4 | csa_tree_add_86_2_n_35);
 assign csa_tree_add_86_2_n_54 = ~(csa_tree_add_86_2_n_27 | csa_tree_add_86_2_n_31);
 assign csa_tree_add_86_2_n_52 = ~(csa_tree_add_86_2_n_25 | csa_tree_add_86_2_n_12);
 assign csa_tree_add_86_2_n_47 = ~(csa_tree_add_86_2_n_4 | csa_tree_add_86_2_n_21);
 assign csa_tree_add_86_2_n_44 = ~(csa_tree_add_86_2_n_3 | csa_tree_add_86_2_n_20);
 assign csa_tree_add_86_2_n_42 = ~(csa_tree_add_86_2_n_3 | csa_tree_add_86_2_n_21);
 assign csa_tree_add_86_2_n_41 = ~(csa_tree_add_86_2_n_18 | ~{in5[1]});
 assign csa_tree_add_86_2_n_37 = ~n_1349;
 assign csa_tree_add_86_2_n_35 = ~n_1347;
 assign csa_tree_add_86_2_n_34 = ~n_1330;
 assign csa_tree_add_86_2_n_33 = ~n_1346;
 assign csa_tree_add_86_2_n_31 = ~n_1344;
 assign csa_tree_add_86_2_n_30 = ~n_1325;
 assign csa_tree_add_86_2_n_23 = ~n_1335;
 assign csa_tree_add_86_2_n_21 = ~n_1497;
 assign csa_tree_add_86_2_n_20 = ~n_1348;
 assign csa_tree_add_86_2_n_19 = ~n_1327;
 assign csa_tree_add_86_2_n_18 = ~n_1495;
 assign csa_tree_add_86_2_n_17 = ~n_1329;
 assign csa_tree_add_86_2_n_16 = ~n_1333;
 assign csa_tree_add_86_2_n_15 = ~n_1328;
 assign csa_tree_add_86_2_n_14 = ~n_1326;
 assign csa_tree_add_86_2_n_12 = ~n_1496;
 assign csa_tree_add_86_2_n_11 = ~n_1350;
 assign csa_tree_add_86_2_n_10 = ~n_1332;
 assign csa_tree_add_86_2_n_9 = ~n_1331;
 assign csa_tree_add_86_2_n_8 = ~n_1334;
 assign csa_tree_add_92_2_groupi_n_282 = ((csa_tree_add_92_2_groupi_n_280 & csa_tree_add_92_2_groupi_n_89)
    | ((csa_tree_add_92_2_groupi_n_89 & csa_tree_add_92_2_groupi_n_65) | (csa_tree_add_92_2_groupi_n_65 &
    csa_tree_add_92_2_groupi_n_280)));
 assign n_1408 = (csa_tree_add_92_2_groupi_n_89 ^ (csa_tree_add_92_2_groupi_n_65 ^ csa_tree_add_92_2_groupi_n_280));
 assign csa_tree_add_92_2_groupi_n_280 = ((csa_tree_add_92_2_groupi_n_278 & csa_tree_add_92_2_groupi_n_81)
    | ((csa_tree_add_92_2_groupi_n_81 & csa_tree_add_92_2_groupi_n_90) | (csa_tree_add_92_2_groupi_n_90 &
    csa_tree_add_92_2_groupi_n_278)));
 assign n_1409 = (csa_tree_add_92_2_groupi_n_81 ^ (csa_tree_add_92_2_groupi_n_90 ^ csa_tree_add_92_2_groupi_n_278));
 assign csa_tree_add_92_2_groupi_n_278 = ((csa_tree_add_92_2_groupi_n_276 & csa_tree_add_92_2_groupi_n_91)
    | ((csa_tree_add_92_2_groupi_n_91 & csa_tree_add_92_2_groupi_n_82) | (csa_tree_add_92_2_groupi_n_82 &
    csa_tree_add_92_2_groupi_n_276)));
 assign n_1410 = (csa_tree_add_92_2_groupi_n_91 ^ (csa_tree_add_92_2_groupi_n_82 ^ csa_tree_add_92_2_groupi_n_276));
 assign csa_tree_add_92_2_groupi_n_226 = ((csa_tree_add_92_2_groupi_n_199 & n_1399) | ((n_1399 & csa_tree_add_92_2_groupi_n_208)
    | (csa_tree_add_92_2_groupi_n_208 & csa_tree_add_92_2_groupi_n_199)));
 assign csa_tree_add_92_2_groupi_n_227 = (n_1399 ^ (csa_tree_add_92_2_groupi_n_208 ^ csa_tree_add_92_2_groupi_n_199));
 assign csa_tree_add_92_2_groupi_n_220 = ((csa_tree_add_92_2_groupi_n_198 & csa_tree_add_92_2_groupi_n_195)
    | ((csa_tree_add_92_2_groupi_n_195 & n_1367) | (n_1367 & csa_tree_add_92_2_groupi_n_198)));
 assign csa_tree_add_92_2_groupi_n_221 = (csa_tree_add_92_2_groupi_n_195 ^ (n_1367 ^ csa_tree_add_92_2_groupi_n_198));
 assign csa_tree_add_92_2_groupi_n_210 = ((csa_tree_add_92_2_groupi_n_189 & csa_tree_add_92_2_groupi_n_194)
    | ((csa_tree_add_92_2_groupi_n_194 & n_1397) | (n_1397 & csa_tree_add_92_2_groupi_n_189)));
 assign csa_tree_add_92_2_groupi_n_211 = (csa_tree_add_92_2_groupi_n_194 ^ (n_1397 ^ csa_tree_add_92_2_groupi_n_189));
 assign csa_tree_add_92_2_groupi_n_206 = ((csa_tree_add_92_2_groupi_n_196 & csa_tree_add_92_2_groupi_n_166)
    | ((csa_tree_add_92_2_groupi_n_166 & csa_tree_add_92_2_groupi_n_187) | (csa_tree_add_92_2_groupi_n_187
    & csa_tree_add_92_2_groupi_n_196)));
 assign csa_tree_add_92_2_groupi_n_207 = (csa_tree_add_92_2_groupi_n_166 ^ (csa_tree_add_92_2_groupi_n_187
    ^ csa_tree_add_92_2_groupi_n_196));
 assign csa_tree_add_92_2_groupi_n_204 = ((csa_tree_add_92_2_groupi_n_188 & csa_tree_add_92_2_groupi_n_165)
    | ((csa_tree_add_92_2_groupi_n_165 & n_1396) | (n_1396 & csa_tree_add_92_2_groupi_n_188)));
 assign csa_tree_add_92_2_groupi_n_205 = (csa_tree_add_92_2_groupi_n_165 ^ (n_1396 ^ csa_tree_add_92_2_groupi_n_188));
 assign csa_tree_add_92_2_groupi_n_202 = ((csa_tree_add_92_2_groupi_n_185 & n_1402) | ((n_1402 & n_1372)
    | (n_1372 & csa_tree_add_92_2_groupi_n_185)));
 assign csa_tree_add_92_2_groupi_n_203 = (n_1402 ^ (n_1372 ^ csa_tree_add_92_2_groupi_n_185));
 assign csa_tree_add_92_2_groupi_n_196 = ((csa_tree_add_92_2_groupi_n_184 & csa_tree_add_92_2_groupi_n_161)
    | ((csa_tree_add_92_2_groupi_n_161 & csa_tree_add_92_2_groupi_n_167) | (csa_tree_add_92_2_groupi_n_167
    & csa_tree_add_92_2_groupi_n_184)));
 assign csa_tree_add_92_2_groupi_n_197 = (csa_tree_add_92_2_groupi_n_161 ^ (csa_tree_add_92_2_groupi_n_167
    ^ csa_tree_add_92_2_groupi_n_184));
 assign csa_tree_add_92_2_groupi_n_192 = ((csa_tree_add_92_2_groupi_n_171 & n_1403) | ((n_1403 & n_1373)
    | (n_1373 & csa_tree_add_92_2_groupi_n_171)));
 assign csa_tree_add_92_2_groupi_n_193 = (n_1403 ^ (n_1373 ^ csa_tree_add_92_2_groupi_n_171));
 assign csa_tree_add_92_2_groupi_n_186 = ((csa_tree_add_92_2_groupi_n_157 & csa_tree_add_92_2_groupi_n_160)
    | ((csa_tree_add_92_2_groupi_n_160 & csa_tree_add_92_2_groupi_n_137) | (csa_tree_add_92_2_groupi_n_137
    & csa_tree_add_92_2_groupi_n_157)));
 assign csa_tree_add_92_2_groupi_n_187 = (csa_tree_add_92_2_groupi_n_160 ^ (csa_tree_add_92_2_groupi_n_137
    ^ csa_tree_add_92_2_groupi_n_157));
 assign csa_tree_add_92_2_groupi_n_184 = ((csa_tree_add_92_2_groupi_n_170 & csa_tree_add_92_2_groupi_n_138)
    | ((csa_tree_add_92_2_groupi_n_138 & csa_tree_add_92_2_groupi_n_155) | (csa_tree_add_92_2_groupi_n_155
    & csa_tree_add_92_2_groupi_n_170)));
 assign csa_tree_add_92_2_groupi_n_185 = (csa_tree_add_92_2_groupi_n_138 ^ (csa_tree_add_92_2_groupi_n_155
    ^ csa_tree_add_92_2_groupi_n_170));
 assign csa_tree_add_92_2_groupi_n_182 = ((csa_tree_add_92_2_groupi_n_159 & csa_tree_add_92_2_groupi_n_156)
    | ((csa_tree_add_92_2_groupi_n_156 & csa_tree_add_92_2_groupi_n_153) | (csa_tree_add_92_2_groupi_n_153
    & csa_tree_add_92_2_groupi_n_159)));
 assign csa_tree_add_92_2_groupi_n_183 = (csa_tree_add_92_2_groupi_n_156 ^ (csa_tree_add_92_2_groupi_n_153
    ^ csa_tree_add_92_2_groupi_n_159));
 assign csa_tree_add_92_2_groupi_n_176 = ((csa_tree_add_92_2_groupi_n_164 & n_1395) | ((n_1395 & n_1364)
    | (n_1364 & csa_tree_add_92_2_groupi_n_164)));
 assign csa_tree_add_92_2_groupi_n_177 = (n_1395 ^ (n_1364 ^ csa_tree_add_92_2_groupi_n_164));
 assign csa_tree_add_92_2_groupi_n_174 = ((csa_tree_add_92_2_groupi_n_151 & n_1404) | ((n_1404 & n_1374)
    | (n_1374 & csa_tree_add_92_2_groupi_n_151)));
 assign csa_tree_add_92_2_groupi_n_175 = (n_1404 ^ (n_1374 ^ csa_tree_add_92_2_groupi_n_151));
 assign csa_tree_add_92_2_groupi_n_170 = ((csa_tree_add_92_2_groupi_n_150 & csa_tree_add_92_2_groupi_n_123)
    | ((csa_tree_add_92_2_groupi_n_123 & csa_tree_add_92_2_groupi_n_139) | (csa_tree_add_92_2_groupi_n_139
    & csa_tree_add_92_2_groupi_n_150)));
 assign csa_tree_add_92_2_groupi_n_171 = (csa_tree_add_92_2_groupi_n_123 ^ (csa_tree_add_92_2_groupi_n_139
    ^ csa_tree_add_92_2_groupi_n_150));
 assign csa_tree_add_92_2_groupi_n_168 = ((csa_tree_add_92_2_groupi_n_152 & csa_tree_add_92_2_groupi_n_128)
    | ((csa_tree_add_92_2_groupi_n_128 & csa_tree_add_92_2_groupi_n_105) | (csa_tree_add_92_2_groupi_n_105
    & csa_tree_add_92_2_groupi_n_152)));
 assign csa_tree_add_92_2_groupi_n_169 = (csa_tree_add_92_2_groupi_n_128 ^ (csa_tree_add_92_2_groupi_n_105
    ^ csa_tree_add_92_2_groupi_n_152));
 assign csa_tree_add_92_2_groupi_n_166 = ((csa_tree_add_92_2_groupi_n_154 & csa_tree_add_92_2_groupi_n_133)
    | ((csa_tree_add_92_2_groupi_n_133 & csa_tree_add_92_2_groupi_n_113) | (csa_tree_add_92_2_groupi_n_113
    & csa_tree_add_92_2_groupi_n_154)));
 assign csa_tree_add_92_2_groupi_n_167 = (csa_tree_add_92_2_groupi_n_133 ^ (csa_tree_add_92_2_groupi_n_113
    ^ csa_tree_add_92_2_groupi_n_154));
 assign csa_tree_add_92_2_groupi_n_160 = ((csa_tree_add_92_2_groupi_n_126 & csa_tree_add_92_2_groupi_n_130)
    | ((csa_tree_add_92_2_groupi_n_130 & csa_tree_add_92_2_groupi_n_12) | (csa_tree_add_92_2_groupi_n_12
    & csa_tree_add_92_2_groupi_n_126)));
 assign csa_tree_add_92_2_groupi_n_161 = (csa_tree_add_92_2_groupi_n_130 ^ (csa_tree_add_92_2_groupi_n_12
    ^ csa_tree_add_92_2_groupi_n_126));
 assign csa_tree_add_92_2_groupi_n_158 = ((csa_tree_add_92_2_groupi_n_136 & csa_tree_add_92_2_groupi_n_129)
    | ((csa_tree_add_92_2_groupi_n_129 & csa_tree_add_92_2_groupi_n_115) | (csa_tree_add_92_2_groupi_n_115
    & csa_tree_add_92_2_groupi_n_136)));
 assign csa_tree_add_92_2_groupi_n_159 = (csa_tree_add_92_2_groupi_n_129 ^ (csa_tree_add_92_2_groupi_n_115
    ^ csa_tree_add_92_2_groupi_n_136));
 assign csa_tree_add_92_2_groupi_n_156 = ((csa_tree_add_92_2_groupi_n_125 & csa_tree_add_92_2_groupi_n_132)
    | ((csa_tree_add_92_2_groupi_n_132 & csa_tree_add_92_2_groupi_n_111) | (csa_tree_add_92_2_groupi_n_111
    & csa_tree_add_92_2_groupi_n_125)));
 assign csa_tree_add_92_2_groupi_n_157 = (csa_tree_add_92_2_groupi_n_132 ^ (csa_tree_add_92_2_groupi_n_111
    ^ csa_tree_add_92_2_groupi_n_125));
 assign csa_tree_add_92_2_groupi_n_154 = ((csa_tree_add_92_2_groupi_n_131 & csa_tree_add_92_2_groupi_n_127)
    | ((csa_tree_add_92_2_groupi_n_127 & csa_tree_add_92_2_groupi_n_122) | (csa_tree_add_92_2_groupi_n_122
    & csa_tree_add_92_2_groupi_n_131)));
 assign csa_tree_add_92_2_groupi_n_155 = (csa_tree_add_92_2_groupi_n_127 ^ (csa_tree_add_92_2_groupi_n_122
    ^ csa_tree_add_92_2_groupi_n_131));
 assign csa_tree_add_92_2_groupi_n_152 = ((csa_tree_add_92_2_groupi_n_124 & csa_tree_add_92_2_groupi_n_6)
    | ((csa_tree_add_92_2_groupi_n_6 & csa_tree_add_92_2_groupi_n_110) | (csa_tree_add_92_2_groupi_n_110
    & csa_tree_add_92_2_groupi_n_124)));
 assign csa_tree_add_92_2_groupi_n_153 = (csa_tree_add_92_2_groupi_n_6 ^ (csa_tree_add_92_2_groupi_n_110
    ^ csa_tree_add_92_2_groupi_n_124));
 assign csa_tree_add_92_2_groupi_n_150 = ((csa_tree_add_92_2_groupi_n_116 & csa_tree_add_92_2_groupi_n_119)
    | ((csa_tree_add_92_2_groupi_n_119 & csa_tree_add_92_2_groupi_n_24) | (csa_tree_add_92_2_groupi_n_24
    & csa_tree_add_92_2_groupi_n_116)));
 assign csa_tree_add_92_2_groupi_n_151 = (csa_tree_add_92_2_groupi_n_119 ^ (csa_tree_add_92_2_groupi_n_24
    ^ csa_tree_add_92_2_groupi_n_116));
 assign csa_tree_add_92_2_groupi_n_148 = ((csa_tree_add_92_2_groupi_n_117 & n_1405) | ((n_1405 & csa_tree_add_92_2_groupi_n_98)
    | (csa_tree_add_92_2_groupi_n_98 & csa_tree_add_92_2_groupi_n_117)));
 assign csa_tree_add_92_2_groupi_n_149 = (n_1405 ^ (csa_tree_add_92_2_groupi_n_98 ^ csa_tree_add_92_2_groupi_n_117));
 assign csa_tree_add_92_2_groupi_n_146 = ((csa_tree_add_92_2_groupi_n_103 & csa_tree_add_92_2_groupi_n_104)
    | ((csa_tree_add_92_2_groupi_n_104 & csa_tree_add_92_2_groupi_n_121) | (csa_tree_add_92_2_groupi_n_121
    & csa_tree_add_92_2_groupi_n_103)));
 assign csa_tree_add_92_2_groupi_n_147 = (csa_tree_add_92_2_groupi_n_104 ^ (csa_tree_add_92_2_groupi_n_121
    ^ csa_tree_add_92_2_groupi_n_103));
 assign csa_tree_add_92_2_groupi_n_144 = ((csa_tree_add_92_2_groupi_n_102 & csa_tree_add_92_2_groupi_n_107)
    | ((csa_tree_add_92_2_groupi_n_107 & csa_tree_add_92_2_groupi_n_7) | (csa_tree_add_92_2_groupi_n_7 &
    csa_tree_add_92_2_groupi_n_102)));
 assign csa_tree_add_92_2_groupi_n_145 = (csa_tree_add_92_2_groupi_n_107 ^ (csa_tree_add_92_2_groupi_n_7
    ^ csa_tree_add_92_2_groupi_n_102));
 assign csa_tree_add_92_2_groupi_n_140 = ((csa_tree_add_92_2_groupi_n_114 & csa_tree_add_92_2_groupi_n_46)
    | ((csa_tree_add_92_2_groupi_n_46 & csa_tree_add_92_2_groupi_n_96) | (csa_tree_add_92_2_groupi_n_96 &
    csa_tree_add_92_2_groupi_n_114)));
 assign csa_tree_add_92_2_groupi_n_141 = (csa_tree_add_92_2_groupi_n_46 ^ (csa_tree_add_92_2_groupi_n_96
    ^ csa_tree_add_92_2_groupi_n_114));
 assign csa_tree_add_92_2_groupi_n_138 = ((csa_tree_add_92_2_groupi_n_118 & csa_tree_add_92_2_groupi_n_35)
    | ((csa_tree_add_92_2_groupi_n_35 & csa_tree_add_92_2_groupi_n_8) | (csa_tree_add_92_2_groupi_n_8 & csa_tree_add_92_2_groupi_n_118)));
 assign csa_tree_add_92_2_groupi_n_139 = (csa_tree_add_92_2_groupi_n_35 ^ (csa_tree_add_92_2_groupi_n_8
    ^ csa_tree_add_92_2_groupi_n_118));
 assign csa_tree_add_92_2_groupi_n_136 = ((csa_tree_add_92_2_groupi_n_112 & csa_tree_add_92_2_groupi_n_4)
    | ((csa_tree_add_92_2_groupi_n_4 & csa_tree_add_92_2_groupi_n_38) | (csa_tree_add_92_2_groupi_n_38 &
    csa_tree_add_92_2_groupi_n_112)));
 assign csa_tree_add_92_2_groupi_n_137 = (csa_tree_add_92_2_groupi_n_4 ^ (csa_tree_add_92_2_groupi_n_38
    ^ csa_tree_add_92_2_groupi_n_112));
 assign csa_tree_add_92_2_groupi_n_132 = ((csa_tree_add_92_2_groupi_n_55 & csa_tree_add_92_2_groupi_n_20)
    | ((csa_tree_add_92_2_groupi_n_20 & csa_tree_add_92_2_groupi_n_39) | (csa_tree_add_92_2_groupi_n_39 &
    csa_tree_add_92_2_groupi_n_55)));
 assign csa_tree_add_92_2_groupi_n_133 = (csa_tree_add_92_2_groupi_n_20 ^ (csa_tree_add_92_2_groupi_n_39
    ^ csa_tree_add_92_2_groupi_n_55));
 assign csa_tree_add_92_2_groupi_n_130 = ((csa_tree_add_92_2_groupi_n_52 & csa_tree_add_92_2_groupi_n_22)
    | ((csa_tree_add_92_2_groupi_n_22 & csa_tree_add_92_2_groupi_n_49) | (csa_tree_add_92_2_groupi_n_49 &
    csa_tree_add_92_2_groupi_n_52)));
 assign csa_tree_add_92_2_groupi_n_131 = (csa_tree_add_92_2_groupi_n_22 ^ (csa_tree_add_92_2_groupi_n_49
    ^ csa_tree_add_92_2_groupi_n_52));
 assign csa_tree_add_92_2_groupi_n_128 = ((csa_tree_add_92_2_groupi_n_50 & csa_tree_add_92_2_groupi_n_45)
    | ((csa_tree_add_92_2_groupi_n_45 & csa_tree_add_92_2_groupi_n_26) | (csa_tree_add_92_2_groupi_n_26 &
    csa_tree_add_92_2_groupi_n_50)));
 assign csa_tree_add_92_2_groupi_n_129 = (csa_tree_add_92_2_groupi_n_45 ^ (csa_tree_add_92_2_groupi_n_26
    ^ csa_tree_add_92_2_groupi_n_50));
 assign csa_tree_add_92_2_groupi_n_126 = ((csa_tree_add_92_2_groupi_n_58 & csa_tree_add_92_2_groupi_n_23)
    | ((csa_tree_add_92_2_groupi_n_23 & csa_tree_add_92_2_groupi_n_1) | (csa_tree_add_92_2_groupi_n_1 & csa_tree_add_92_2_groupi_n_58)));
 assign csa_tree_add_92_2_groupi_n_127 = (csa_tree_add_92_2_groupi_n_23 ^ (csa_tree_add_92_2_groupi_n_1
    ^ csa_tree_add_92_2_groupi_n_58));
 assign csa_tree_add_92_2_groupi_n_124 = ((csa_tree_add_92_2_groupi_n_61 & csa_tree_add_92_2_groupi_n_40)
    | ((csa_tree_add_92_2_groupi_n_40 & csa_tree_add_92_2_groupi_n_2) | (csa_tree_add_92_2_groupi_n_2 & csa_tree_add_92_2_groupi_n_61)));
 assign csa_tree_add_92_2_groupi_n_125 = (csa_tree_add_92_2_groupi_n_40 ^ (csa_tree_add_92_2_groupi_n_2
    ^ csa_tree_add_92_2_groupi_n_61));
 assign csa_tree_add_92_2_groupi_n_122 = ((csa_tree_add_92_2_groupi_n_54 & csa_tree_add_92_2_groupi_n_19)
    | ((csa_tree_add_92_2_groupi_n_19 & csa_tree_add_92_2_groupi_n_13) | (csa_tree_add_92_2_groupi_n_13 &
    csa_tree_add_92_2_groupi_n_54)));
 assign csa_tree_add_92_2_groupi_n_123 = (csa_tree_add_92_2_groupi_n_19 ^ (csa_tree_add_92_2_groupi_n_13
    ^ csa_tree_add_92_2_groupi_n_54));
 assign csa_tree_add_92_2_groupi_n_120 = ((csa_tree_add_92_2_groupi_n_95 & csa_tree_add_92_2_groupi_n_47)
    | ((csa_tree_add_92_2_groupi_n_47 & csa_tree_add_92_2_groupi_n_25) | (csa_tree_add_92_2_groupi_n_25 &
    csa_tree_add_92_2_groupi_n_95)));
 assign csa_tree_add_92_2_groupi_n_121 = (csa_tree_add_92_2_groupi_n_47 ^ (csa_tree_add_92_2_groupi_n_25
    ^ csa_tree_add_92_2_groupi_n_95));
 assign csa_tree_add_92_2_groupi_n_118 = ((csa_tree_add_92_2_groupi_n_63 & csa_tree_add_92_2_groupi_n_3)
    | ((csa_tree_add_92_2_groupi_n_3 & csa_tree_add_92_2_groupi_n_21) | (csa_tree_add_92_2_groupi_n_21 &
    csa_tree_add_92_2_groupi_n_63)));
 assign csa_tree_add_92_2_groupi_n_119 = (csa_tree_add_92_2_groupi_n_3 ^ (csa_tree_add_92_2_groupi_n_21
    ^ csa_tree_add_92_2_groupi_n_63));
 assign csa_tree_add_92_2_groupi_n_116 = ((csa_tree_add_92_2_groupi_n_28 & csa_tree_add_92_2_groupi_n_27)
    | ((csa_tree_add_92_2_groupi_n_27 & csa_tree_add_92_2_groupi_n_18) | (csa_tree_add_92_2_groupi_n_18 &
    csa_tree_add_92_2_groupi_n_28)));
 assign csa_tree_add_92_2_groupi_n_117 = (csa_tree_add_92_2_groupi_n_27 ^ (csa_tree_add_92_2_groupi_n_18
    ^ csa_tree_add_92_2_groupi_n_28));
 assign csa_tree_add_92_2_groupi_n_114 = ((csa_tree_add_92_2_groupi_n_57 & csa_tree_add_92_2_groupi_n_48)
    | ((csa_tree_add_92_2_groupi_n_48 & csa_tree_add_92_2_groupi_n_33) | (csa_tree_add_92_2_groupi_n_33 &
    csa_tree_add_92_2_groupi_n_57)));
 assign csa_tree_add_92_2_groupi_n_115 = (csa_tree_add_92_2_groupi_n_48 ^ (csa_tree_add_92_2_groupi_n_33
    ^ csa_tree_add_92_2_groupi_n_57));
 assign csa_tree_add_92_2_groupi_n_112 = ((csa_tree_add_92_2_groupi_n_51 & csa_tree_add_92_2_groupi_n_17)
    | ((csa_tree_add_92_2_groupi_n_17 & csa_tree_add_92_2_groupi_n_15) | (csa_tree_add_92_2_groupi_n_15 &
    csa_tree_add_92_2_groupi_n_51)));
 assign csa_tree_add_92_2_groupi_n_113 = (csa_tree_add_92_2_groupi_n_17 ^ (csa_tree_add_92_2_groupi_n_15
    ^ csa_tree_add_92_2_groupi_n_51));
 assign csa_tree_add_92_2_groupi_n_110 = ((csa_tree_add_92_2_groupi_n_59 & csa_tree_add_92_2_groupi_n_43)
    | ((csa_tree_add_92_2_groupi_n_43 & csa_tree_add_92_2_groupi_n_14) | (csa_tree_add_92_2_groupi_n_14 &
    csa_tree_add_92_2_groupi_n_59)));
 assign csa_tree_add_92_2_groupi_n_111 = (csa_tree_add_92_2_groupi_n_43 ^ (csa_tree_add_92_2_groupi_n_14
    ^ csa_tree_add_92_2_groupi_n_59));
 assign csa_tree_add_92_2_groupi_n_108 = ((csa_tree_add_92_2_groupi_n_29 & csa_tree_add_92_2_groupi_n_9)
    | ((csa_tree_add_92_2_groupi_n_9 & csa_tree_add_92_2_groupi_n_10) | (csa_tree_add_92_2_groupi_n_10 &
    csa_tree_add_92_2_groupi_n_29)));
 assign csa_tree_add_92_2_groupi_n_109 = (csa_tree_add_92_2_groupi_n_9 ^ (csa_tree_add_92_2_groupi_n_10
    ^ csa_tree_add_92_2_groupi_n_29));
 assign csa_tree_add_92_2_groupi_n_106 = ((csa_tree_add_92_2_groupi_n_56 & csa_tree_add_92_2_groupi_n_36)
    | ((csa_tree_add_92_2_groupi_n_36 & csa_tree_add_92_2_groupi_n_37) | (csa_tree_add_92_2_groupi_n_37 &
    csa_tree_add_92_2_groupi_n_56)));
 assign csa_tree_add_92_2_groupi_n_107 = (csa_tree_add_92_2_groupi_n_36 ^ (csa_tree_add_92_2_groupi_n_37
    ^ csa_tree_add_92_2_groupi_n_56));
 assign csa_tree_add_92_2_groupi_n_104 = ((csa_tree_add_92_2_groupi_n_53 & csa_tree_add_92_2_groupi_n_34)
    | ((csa_tree_add_92_2_groupi_n_34 & csa_tree_add_92_2_groupi_n_5) | (csa_tree_add_92_2_groupi_n_5 & csa_tree_add_92_2_groupi_n_53)));
 assign csa_tree_add_92_2_groupi_n_105 = (csa_tree_add_92_2_groupi_n_34 ^ (csa_tree_add_92_2_groupi_n_5
    ^ csa_tree_add_92_2_groupi_n_53));
 assign csa_tree_add_92_2_groupi_n_102 = ((csa_tree_add_92_2_groupi_n_62 & csa_tree_add_92_2_groupi_n_0)
    | ((csa_tree_add_92_2_groupi_n_0 & csa_tree_add_92_2_groupi_n_16) | (csa_tree_add_92_2_groupi_n_16 &
    csa_tree_add_92_2_groupi_n_62)));
 assign csa_tree_add_92_2_groupi_n_103 = (csa_tree_add_92_2_groupi_n_0 ^ (csa_tree_add_92_2_groupi_n_16
    ^ csa_tree_add_92_2_groupi_n_62));
 assign csa_tree_add_92_2_groupi_n_98 = ((csa_tree_add_92_2_groupi_n_60 & n_1406) | ((n_1406 & csa_tree_add_92_2_groupi_n_41)
    | (csa_tree_add_92_2_groupi_n_41 & csa_tree_add_92_2_groupi_n_60)));
 assign csa_tree_add_92_2_groupi_n_99 = (n_1406 ^ (csa_tree_add_92_2_groupi_n_41 ^ csa_tree_add_92_2_groupi_n_60));
 assign csa_tree_add_92_2_groupi_n_95 = (csa_tree_add_92_2_groupi_n_64 & csa_tree_add_92_2_groupi_n_30);
 assign csa_tree_add_92_2_groupi_n_96 = (csa_tree_add_92_2_groupi_n_64 ^ csa_tree_add_92_2_groupi_n_30);
 assign csa_tree_add_92_2_groupi_n_93 = (n_1385 & n_1354);
 assign csa_tree_add_92_2_groupi_n_94 = (n_1385 ^ n_1354);
 assign csa_tree_add_92_2_groupi_n_87 = (n_1388 & n_1357);
 assign csa_tree_add_92_2_groupi_n_88 = (n_1388 ^ n_1357);
 assign csa_tree_add_92_2_groupi_n_85 = (n_1390 & n_1359);
 assign csa_tree_add_92_2_groupi_n_86 = (n_1390 ^ n_1359);
 assign csa_tree_add_92_2_groupi_n_83 = (n_1387 & n_1356);
 assign csa_tree_add_92_2_groupi_n_84 = (n_1387 ^ n_1356);
 assign csa_tree_add_92_2_groupi_n_79 = (n_1386 & n_1355);
 assign csa_tree_add_92_2_groupi_n_80 = (n_1386 ^ n_1355);
 assign csa_tree_add_92_2_groupi_n_77 = (n_1394 & n_1363);
 assign csa_tree_add_92_2_groupi_n_78 = (n_1394 ^ n_1363);
 assign csa_tree_add_92_2_groupi_n_73 = (n_1392 & n_1361);
 assign csa_tree_add_92_2_groupi_n_74 = (n_1392 ^ n_1361);
 assign csa_tree_add_92_2_groupi_n_71 = (n_1391 & n_1360);
 assign csa_tree_add_92_2_groupi_n_72 = (n_1391 ^ n_1360);
 assign csa_tree_add_92_2_groupi_n_69 = (n_1393 & n_1362);
 assign csa_tree_add_92_2_groupi_n_70 = (n_1393 ^ n_1362);
 assign csa_tree_add_92_2_groupi_n_67 = (n_1389 & n_1358);
 assign csa_tree_add_92_2_groupi_n_68 = (n_1389 ^ n_1358);
 assign csa_tree_add_92_2_groupi_n_66 = ~(n_1379 ^ n_1351);
 assign csa_tree_add_92_2_groupi_n_64 = ({in7[2]} & {in8[7]});
 assign csa_tree_add_92_2_groupi_n_63 = ({in7[3]} & {in8[0]});
 assign csa_tree_add_92_2_groupi_n_62 = ({in7[7]} & {in8[3]});
 assign csa_tree_add_92_2_groupi_n_61 = ({in7[6]} & {in8[1]});
 assign csa_tree_add_92_2_groupi_n_60 = ({in7[1]} & {in8[0]});
 assign csa_tree_add_92_2_groupi_n_59 = ({in7[4]} & {in8[3]});
 assign csa_tree_add_92_2_groupi_n_58 = ({in7[4]} & {in8[1]});
 assign csa_tree_add_92_2_groupi_n_57 = ({in7[3]} & {in8[5]});
 assign csa_tree_add_92_2_groupi_n_56 = ({in7[5]} & {in8[6]});
 assign csa_tree_add_92_2_groupi_n_55 = ({in7[5]} & {in8[1]});
 assign csa_tree_add_92_2_groupi_n_54 = ({in7[1]} & {in8[3]});
 assign csa_tree_add_92_2_groupi_n_53 = ({in7[7]} & {in8[2]});
 assign csa_tree_add_92_2_groupi_n_52 = ({in7[2]} & {in8[3]});
 assign csa_tree_add_92_2_groupi_n_51 = ({in7[2]} & {in8[4]});
 assign csa_tree_add_92_2_groupi_n_50 = ({in7[6]} & {in8[2]});
 assign csa_tree_add_92_2_groupi_n_49 = ({in7[0]} & {in8[5]});
 assign csa_tree_add_92_2_groupi_n_48 = ({in7[7]} & {in8[1]});
 assign csa_tree_add_92_2_groupi_n_47 = ({in7[6]} & {in8[4]});
 assign csa_tree_add_92_2_groupi_n_46 = ({in7[6]} & {in8[3]});
 assign csa_tree_add_92_2_groupi_n_45 = ({in7[5]} & {in8[3]});
 assign csa_tree_add_92_2_groupi_n_43 = ({in7[3]} & {in8[4]});
 assign csa_tree_add_92_2_groupi_n_42 = ({in7[7]} & {in8[6]});
 assign csa_tree_add_92_2_groupi_n_41 = ({in7[0]} & {in8[1]});
 assign csa_tree_add_92_2_groupi_n_40 = ({in7[7]} & {in8[0]});
 assign csa_tree_add_92_2_groupi_n_39 = ({in7[3]} & {in8[3]});
 assign csa_tree_add_92_2_groupi_n_38 = ({in7[1]} & {in8[6]});
 assign csa_tree_add_92_2_groupi_n_37 = ({in7[4]} & {in8[7]});
 assign csa_tree_add_92_2_groupi_n_36 = ({in7[7]} & {in8[4]});
 assign csa_tree_add_92_2_groupi_n_35 = ({in7[3]} & {in8[1]});
 assign csa_tree_add_92_2_groupi_n_34 = ({in7[5]} & {in8[4]});
 assign csa_tree_add_92_2_groupi_n_33 = ({in7[1]} & {in8[7]});
 assign csa_tree_add_92_2_groupi_n_32 = ~(n_1380 & n_1352);
 assign csa_tree_add_92_2_groupi_n_31 = ({in7[0]} & {in8[0]});
 assign csa_tree_add_92_2_groupi_n_30 = ({in7[3]} & {in8[6]});
 assign csa_tree_add_92_2_groupi_n_29 = ({in7[7]} & {in8[5]});
 assign csa_tree_add_92_2_groupi_n_28 = ({in7[1]} & {in8[1]});
 assign csa_tree_add_92_2_groupi_n_27 = ({in7[2]} & {in8[0]});
 assign csa_tree_add_92_2_groupi_n_26 = ({in7[4]} & {in8[4]});
 assign csa_tree_add_92_2_groupi_n_25 = ({in7[5]} & {in8[5]});
 assign csa_tree_add_92_2_groupi_n_24 = ({in7[2]} & {in8[1]});
 assign csa_tree_add_92_2_groupi_n_23 = ({in7[5]} & {in8[0]});
 assign csa_tree_add_92_2_groupi_n_22 = ({in7[1]} & {in8[4]});
 assign csa_tree_add_92_2_groupi_n_21 = ({in7[0]} & {in8[3]});
 assign csa_tree_add_92_2_groupi_n_20 = ({in7[4]} & {in8[2]});
 assign csa_tree_add_92_2_groupi_n_19 = ({in7[4]} & {in8[0]});
 assign csa_tree_add_92_2_groupi_n_18 = ({in7[0]} & {in8[2]});
 assign csa_tree_add_92_2_groupi_n_17 = ({in7[6]} & {in8[0]});
 assign csa_tree_add_92_2_groupi_n_16 = ({in7[3]} & {in8[7]});
 assign csa_tree_add_92_2_groupi_n_15 = ({in7[0]} & {in8[6]});
 assign csa_tree_add_92_2_groupi_n_14 = ({in7[2]} & {in8[5]});
 assign csa_tree_add_92_2_groupi_n_13 = ({in7[0]} & {in8[4]});
 assign csa_tree_add_92_2_groupi_n_12 = ({in7[1]} & {in8[5]});
 assign csa_tree_add_92_2_groupi_n_11 = ({in7[6]} & {in8[7]});
 assign csa_tree_add_92_2_groupi_n_10 = ({in7[5]} & {in8[7]});
 assign csa_tree_add_92_2_groupi_n_9 = ({in7[6]} & {in8[6]});
 assign csa_tree_add_92_2_groupi_n_8 = ({in7[2]} & {in8[2]});
 assign csa_tree_add_92_2_groupi_n_7 = ({in7[6]} & {in8[5]});
 assign csa_tree_add_92_2_groupi_n_6 = ({in7[2]} & {in8[6]});
 assign csa_tree_add_92_2_groupi_n_5 = ({in7[4]} & {in8[5]});
 assign csa_tree_add_92_2_groupi_n_4 = ({in7[5]} & {in8[2]});
 assign csa_tree_add_92_2_groupi_n_3 = ({in7[1]} & {in8[2]});
 assign csa_tree_add_92_2_groupi_n_2 = ({in7[0]} & {in8[7]});
 assign csa_tree_add_92_2_groupi_n_1 = ({in7[3]} & {in8[2]});
 assign csa_tree_add_92_2_groupi_n_0 = ({in7[4]} & {in8[6]});
 assign n_1448 = ~(csa_tree_add_106_2_groupi_n_1162 ^ csa_tree_add_106_2_groupi_n_1089);
 assign csa_tree_add_106_2_groupi_n_1162 = ((csa_tree_add_106_2_groupi_n_1160 & csa_tree_add_106_2_groupi_n_1076)
    | ((csa_tree_add_106_2_groupi_n_1076 & csa_tree_add_106_2_groupi_n_1079) | (csa_tree_add_106_2_groupi_n_1079
    & csa_tree_add_106_2_groupi_n_1160)));
 assign n_1449 = (csa_tree_add_106_2_groupi_n_1076 ^ (csa_tree_add_106_2_groupi_n_1079 ^ csa_tree_add_106_2_groupi_n_1160));
 assign csa_tree_add_106_2_groupi_n_1160 = ((csa_tree_add_106_2_groupi_n_1158 & csa_tree_add_106_2_groupi_n_1085)
    | ((csa_tree_add_106_2_groupi_n_1085 & csa_tree_add_106_2_groupi_n_1080) | (csa_tree_add_106_2_groupi_n_1080
    & csa_tree_add_106_2_groupi_n_1158)));
 assign n_1450 = (csa_tree_add_106_2_groupi_n_1085 ^ (csa_tree_add_106_2_groupi_n_1080 ^ csa_tree_add_106_2_groupi_n_1158));
 assign csa_tree_add_106_2_groupi_n_1158 = ((csa_tree_add_106_2_groupi_n_1156 & csa_tree_add_106_2_groupi_n_1086)
    | ((csa_tree_add_106_2_groupi_n_1086 & csa_tree_add_106_2_groupi_n_1053) | (csa_tree_add_106_2_groupi_n_1053
    & csa_tree_add_106_2_groupi_n_1156)));
 assign n_1451 = (csa_tree_add_106_2_groupi_n_1086 ^ (csa_tree_add_106_2_groupi_n_1053 ^ csa_tree_add_106_2_groupi_n_1156));
 assign csa_tree_add_106_2_groupi_n_1156 = ((csa_tree_add_106_2_groupi_n_1154 & csa_tree_add_106_2_groupi_n_1057)
    | ((csa_tree_add_106_2_groupi_n_1057 & csa_tree_add_106_2_groupi_n_1054) | (csa_tree_add_106_2_groupi_n_1054
    & csa_tree_add_106_2_groupi_n_1154)));
 assign n_1452 = (csa_tree_add_106_2_groupi_n_1057 ^ (csa_tree_add_106_2_groupi_n_1054 ^ csa_tree_add_106_2_groupi_n_1154));
 assign csa_tree_add_106_2_groupi_n_1154 = ((csa_tree_add_106_2_groupi_n_1152 & csa_tree_add_106_2_groupi_n_1058)
    | ((csa_tree_add_106_2_groupi_n_1058 & csa_tree_add_106_2_groupi_n_1087) | (csa_tree_add_106_2_groupi_n_1087
    & csa_tree_add_106_2_groupi_n_1152)));
 assign n_1453 = (csa_tree_add_106_2_groupi_n_1058 ^ (csa_tree_add_106_2_groupi_n_1087 ^ csa_tree_add_106_2_groupi_n_1152));
 assign csa_tree_add_106_2_groupi_n_1152 = ((csa_tree_add_106_2_groupi_n_1150 & csa_tree_add_106_2_groupi_n_1088)
    | ((csa_tree_add_106_2_groupi_n_1088 & csa_tree_add_106_2_groupi_n_1073) | (csa_tree_add_106_2_groupi_n_1073
    & csa_tree_add_106_2_groupi_n_1150)));
 assign n_1454 = (csa_tree_add_106_2_groupi_n_1088 ^ (csa_tree_add_106_2_groupi_n_1073 ^ csa_tree_add_106_2_groupi_n_1150));
 assign csa_tree_add_106_2_groupi_n_1120 = ((csa_tree_add_106_2_groupi_n_1091 & csa_tree_add_106_2_groupi_n_1002)
    | ((csa_tree_add_106_2_groupi_n_1002 & csa_tree_add_106_2_groupi_n_1102) | (csa_tree_add_106_2_groupi_n_1102
    & csa_tree_add_106_2_groupi_n_1091)));
 assign csa_tree_add_106_2_groupi_n_1121 = (csa_tree_add_106_2_groupi_n_1002 ^ (csa_tree_add_106_2_groupi_n_1102
    ^ csa_tree_add_106_2_groupi_n_1091));
 assign csa_tree_add_106_2_groupi_n_1118 = ((csa_tree_add_106_2_groupi_n_1100 & csa_tree_add_106_2_groupi_n_1103)
    | ((csa_tree_add_106_2_groupi_n_1103 & csa_tree_add_106_2_groupi_n_1044) | (csa_tree_add_106_2_groupi_n_1044
    & csa_tree_add_106_2_groupi_n_1100)));
 assign csa_tree_add_106_2_groupi_n_1119 = (csa_tree_add_106_2_groupi_n_1103 ^ (csa_tree_add_106_2_groupi_n_1044
    ^ csa_tree_add_106_2_groupi_n_1100));
 assign csa_tree_add_106_2_groupi_n_1114 = ((csa_tree_add_106_2_groupi_n_1096 & csa_tree_add_106_2_groupi_n_988)
    | ((csa_tree_add_106_2_groupi_n_988 & csa_tree_add_106_2_groupi_n_965) | (csa_tree_add_106_2_groupi_n_965
    & csa_tree_add_106_2_groupi_n_1096)));
 assign csa_tree_add_106_2_groupi_n_1115 = (csa_tree_add_106_2_groupi_n_988 ^ (csa_tree_add_106_2_groupi_n_965
    ^ csa_tree_add_106_2_groupi_n_1096));
 assign csa_tree_add_106_2_groupi_n_1112 = ((csa_tree_add_106_2_groupi_n_1101 & csa_tree_add_106_2_groupi_n_1067)
    | ((csa_tree_add_106_2_groupi_n_1067 & csa_tree_add_106_2_groupi_n_1072) | (csa_tree_add_106_2_groupi_n_1072
    & csa_tree_add_106_2_groupi_n_1101)));
 assign csa_tree_add_106_2_groupi_n_1113 = (csa_tree_add_106_2_groupi_n_1067 ^ (csa_tree_add_106_2_groupi_n_1072
    ^ csa_tree_add_106_2_groupi_n_1101));
 assign csa_tree_add_106_2_groupi_n_1110 = ((csa_tree_add_106_2_groupi_n_1078 & csa_tree_add_106_2_groupi_n_1090)
    | ((csa_tree_add_106_2_groupi_n_1090 & csa_tree_add_106_2_groupi_n_1050) | (csa_tree_add_106_2_groupi_n_1050
    & csa_tree_add_106_2_groupi_n_1078)));
 assign csa_tree_add_106_2_groupi_n_1111 = (csa_tree_add_106_2_groupi_n_1090 ^ (csa_tree_add_106_2_groupi_n_1050
    ^ csa_tree_add_106_2_groupi_n_1078));
 assign csa_tree_add_106_2_groupi_n_1108 = ((csa_tree_add_106_2_groupi_n_1097 & csa_tree_add_106_2_groupi_n_1049)
    | ((csa_tree_add_106_2_groupi_n_1049 & csa_tree_add_106_2_groupi_n_947) | (csa_tree_add_106_2_groupi_n_947
    & csa_tree_add_106_2_groupi_n_1097)));
 assign csa_tree_add_106_2_groupi_n_1109 = (csa_tree_add_106_2_groupi_n_1049 ^ (csa_tree_add_106_2_groupi_n_947
    ^ csa_tree_add_106_2_groupi_n_1097));
 assign csa_tree_add_106_2_groupi_n_1106 = ((csa_tree_add_106_2_groupi_n_1083 & csa_tree_add_106_2_groupi_n_1068)
    | ((csa_tree_add_106_2_groupi_n_1068 & csa_tree_add_106_2_groupi_n_1070) | (csa_tree_add_106_2_groupi_n_1070
    & csa_tree_add_106_2_groupi_n_1083)));
 assign csa_tree_add_106_2_groupi_n_1107 = (csa_tree_add_106_2_groupi_n_1068 ^ (csa_tree_add_106_2_groupi_n_1070
    ^ csa_tree_add_106_2_groupi_n_1083));
 assign csa_tree_add_106_2_groupi_n_1102 = ((csa_tree_add_106_2_groupi_n_1071 & csa_tree_add_106_2_groupi_n_366)
    | ((csa_tree_add_106_2_groupi_n_366 & csa_tree_add_106_2_groupi_n_939) | (csa_tree_add_106_2_groupi_n_939
    & csa_tree_add_106_2_groupi_n_1071)));
 assign csa_tree_add_106_2_groupi_n_1103 = (csa_tree_add_106_2_groupi_n_366 ^ (csa_tree_add_106_2_groupi_n_939
    ^ csa_tree_add_106_2_groupi_n_1071));
 assign csa_tree_add_106_2_groupi_n_1100 = ((csa_tree_add_106_2_groupi_n_1069 & csa_tree_add_106_2_groupi_n_371)
    | ((csa_tree_add_106_2_groupi_n_371 & csa_tree_add_106_2_groupi_n_981) | (csa_tree_add_106_2_groupi_n_981
    & csa_tree_add_106_2_groupi_n_1069)));
 assign csa_tree_add_106_2_groupi_n_1101 = (csa_tree_add_106_2_groupi_n_371 ^ (csa_tree_add_106_2_groupi_n_981
    ^ csa_tree_add_106_2_groupi_n_1069));
 assign csa_tree_add_106_2_groupi_n_1098 = ((csa_tree_add_106_2_groupi_n_1084 & csa_tree_add_106_2_groupi_n_1021)
    | ((csa_tree_add_106_2_groupi_n_1021 & csa_tree_add_106_2_groupi_n_1047) | (csa_tree_add_106_2_groupi_n_1047
    & csa_tree_add_106_2_groupi_n_1084)));
 assign csa_tree_add_106_2_groupi_n_1099 = (csa_tree_add_106_2_groupi_n_1021 ^ (csa_tree_add_106_2_groupi_n_1047
    ^ csa_tree_add_106_2_groupi_n_1084));
 assign csa_tree_add_106_2_groupi_n_1096 = ((csa_tree_add_106_2_groupi_n_1077 & csa_tree_add_106_2_groupi_n_378)
    | ((csa_tree_add_106_2_groupi_n_378 & csa_tree_add_106_2_groupi_n_929) | (csa_tree_add_106_2_groupi_n_929
    & csa_tree_add_106_2_groupi_n_1077)));
 assign csa_tree_add_106_2_groupi_n_1097 = (csa_tree_add_106_2_groupi_n_378 ^ (csa_tree_add_106_2_groupi_n_929
    ^ csa_tree_add_106_2_groupi_n_1077));
 assign csa_tree_add_106_2_groupi_n_1094 = ((csa_tree_add_106_2_groupi_n_1048 & csa_tree_add_106_2_groupi_n_1035)
    | ((csa_tree_add_106_2_groupi_n_1035 & csa_tree_add_106_2_groupi_n_1041) | (csa_tree_add_106_2_groupi_n_1041
    & csa_tree_add_106_2_groupi_n_1048)));
 assign csa_tree_add_106_2_groupi_n_1095 = (csa_tree_add_106_2_groupi_n_1035 ^ (csa_tree_add_106_2_groupi_n_1041
    ^ csa_tree_add_106_2_groupi_n_1048));
 assign csa_tree_add_106_2_groupi_n_1090 = ((csa_tree_add_106_2_groupi_n_1043 & csa_tree_add_106_2_groupi_n_857)
    | ((csa_tree_add_106_2_groupi_n_857 & csa_tree_add_106_2_groupi_n_1031) | (csa_tree_add_106_2_groupi_n_1031
    & csa_tree_add_106_2_groupi_n_1043)));
 assign csa_tree_add_106_2_groupi_n_1091 = (csa_tree_add_106_2_groupi_n_857 ^ (csa_tree_add_106_2_groupi_n_1031
    ^ csa_tree_add_106_2_groupi_n_1043));
 assign csa_tree_add_106_2_groupi_n_1089 = ~(csa_tree_add_106_2_groupi_n_1038 ^ csa_tree_add_106_2_groupi_n_1075);
 assign csa_tree_add_106_2_groupi_n_1083 = ((csa_tree_add_106_2_groupi_n_1025 & csa_tree_add_106_2_groupi_n_369)
    | ((csa_tree_add_106_2_groupi_n_369 & csa_tree_add_106_2_groupi_n_1034) | (csa_tree_add_106_2_groupi_n_1034
    & csa_tree_add_106_2_groupi_n_1025)));
 assign csa_tree_add_106_2_groupi_n_1084 = (csa_tree_add_106_2_groupi_n_369 ^ (csa_tree_add_106_2_groupi_n_1034
    ^ csa_tree_add_106_2_groupi_n_1025));
 assign csa_tree_add_106_2_groupi_n_1081 = ((csa_tree_add_106_2_groupi_n_992 & csa_tree_add_106_2_groupi_n_943)
    | ((csa_tree_add_106_2_groupi_n_943 & csa_tree_add_106_2_groupi_n_1014) | (csa_tree_add_106_2_groupi_n_1014
    & csa_tree_add_106_2_groupi_n_992)));
 assign csa_tree_add_106_2_groupi_n_1082 = (csa_tree_add_106_2_groupi_n_943 ^ (csa_tree_add_106_2_groupi_n_1014
    ^ csa_tree_add_106_2_groupi_n_992));
 assign csa_tree_add_106_2_groupi_n_1079 = ((csa_tree_add_106_2_groupi_n_1022 & csa_tree_add_106_2_groupi_n_1017)
    | ((csa_tree_add_106_2_groupi_n_1017 & csa_tree_add_106_2_groupi_n_963) | (csa_tree_add_106_2_groupi_n_963
    & csa_tree_add_106_2_groupi_n_1022)));
 assign csa_tree_add_106_2_groupi_n_1080 = (csa_tree_add_106_2_groupi_n_1017 ^ (csa_tree_add_106_2_groupi_n_963
    ^ csa_tree_add_106_2_groupi_n_1022));
 assign csa_tree_add_106_2_groupi_n_1077 = ((csa_tree_add_106_2_groupi_n_1030 & csa_tree_add_106_2_groupi_n_377)
    | ((csa_tree_add_106_2_groupi_n_377 & csa_tree_add_106_2_groupi_n_454) | (csa_tree_add_106_2_groupi_n_454
    & csa_tree_add_106_2_groupi_n_1030)));
 assign csa_tree_add_106_2_groupi_n_1078 = (csa_tree_add_106_2_groupi_n_377 ^ (csa_tree_add_106_2_groupi_n_454
    ^ csa_tree_add_106_2_groupi_n_1030));
 assign csa_tree_add_106_2_groupi_n_1075 = ((csa_tree_add_106_2_groupi_n_1016 & csa_tree_add_106_2_groupi_n_1004)
    | ((csa_tree_add_106_2_groupi_n_1004 & csa_tree_add_106_2_groupi_n_973) | (csa_tree_add_106_2_groupi_n_973
    & csa_tree_add_106_2_groupi_n_1016)));
 assign csa_tree_add_106_2_groupi_n_1076 = (csa_tree_add_106_2_groupi_n_1004 ^ (csa_tree_add_106_2_groupi_n_973
    ^ csa_tree_add_106_2_groupi_n_1016));
 assign csa_tree_add_106_2_groupi_n_1071 = ((csa_tree_add_106_2_groupi_n_1028 & csa_tree_add_106_2_groupi_n_451)
    | ((csa_tree_add_106_2_groupi_n_451 & csa_tree_add_106_2_groupi_n_851) | (csa_tree_add_106_2_groupi_n_851
    & csa_tree_add_106_2_groupi_n_1028)));
 assign csa_tree_add_106_2_groupi_n_1072 = (csa_tree_add_106_2_groupi_n_451 ^ (csa_tree_add_106_2_groupi_n_851
    ^ csa_tree_add_106_2_groupi_n_1028));
 assign csa_tree_add_106_2_groupi_n_1069 = ((csa_tree_add_106_2_groupi_n_1024 & csa_tree_add_106_2_groupi_n_446)
    | ((csa_tree_add_106_2_groupi_n_446 & csa_tree_add_106_2_groupi_n_833) | (csa_tree_add_106_2_groupi_n_833
    & csa_tree_add_106_2_groupi_n_1024)));
 assign csa_tree_add_106_2_groupi_n_1070 = (csa_tree_add_106_2_groupi_n_446 ^ (csa_tree_add_106_2_groupi_n_833
    ^ csa_tree_add_106_2_groupi_n_1024));
 assign csa_tree_add_106_2_groupi_n_1067 = ((csa_tree_add_106_2_groupi_n_1029 & csa_tree_add_106_2_groupi_n_368)
    | ((csa_tree_add_106_2_groupi_n_368 & csa_tree_add_106_2_groupi_n_1020) | (csa_tree_add_106_2_groupi_n_1020
    & csa_tree_add_106_2_groupi_n_1029)));
 assign csa_tree_add_106_2_groupi_n_1068 = (csa_tree_add_106_2_groupi_n_368 ^ (csa_tree_add_106_2_groupi_n_1020
    ^ csa_tree_add_106_2_groupi_n_1029));
 assign csa_tree_add_106_2_groupi_n_1063 = ((csa_tree_add_106_2_groupi_n_1042 & csa_tree_add_106_2_groupi_n_367)
    | ((csa_tree_add_106_2_groupi_n_367 & csa_tree_add_106_2_groupi_n_1007) | (csa_tree_add_106_2_groupi_n_1007
    & csa_tree_add_106_2_groupi_n_1042)));
 assign csa_tree_add_106_2_groupi_n_1064 = (csa_tree_add_106_2_groupi_n_367 ^ (csa_tree_add_106_2_groupi_n_1007
    ^ csa_tree_add_106_2_groupi_n_1042));
 assign csa_tree_add_106_2_groupi_n_1057 = ((csa_tree_add_106_2_groupi_n_996 & csa_tree_add_106_2_groupi_n_955)
    | ((csa_tree_add_106_2_groupi_n_955 & csa_tree_add_106_2_groupi_n_989) | (csa_tree_add_106_2_groupi_n_989
    & csa_tree_add_106_2_groupi_n_996)));
 assign csa_tree_add_106_2_groupi_n_1058 = (csa_tree_add_106_2_groupi_n_955 ^ (csa_tree_add_106_2_groupi_n_989
    ^ csa_tree_add_106_2_groupi_n_996));
 assign csa_tree_add_106_2_groupi_n_1053 = ((csa_tree_add_106_2_groupi_n_995 & csa_tree_add_106_2_groupi_n_1027)
    | ((csa_tree_add_106_2_groupi_n_1027 & csa_tree_add_106_2_groupi_n_954) | (csa_tree_add_106_2_groupi_n_954
    & csa_tree_add_106_2_groupi_n_995)));
 assign csa_tree_add_106_2_groupi_n_1054 = (csa_tree_add_106_2_groupi_n_1027 ^ (csa_tree_add_106_2_groupi_n_954
    ^ csa_tree_add_106_2_groupi_n_995));
 assign csa_tree_add_106_2_groupi_n_1051 = ((csa_tree_add_106_2_groupi_n_987 & csa_tree_add_106_2_groupi_n_1015)
    | ((csa_tree_add_106_2_groupi_n_1015 & csa_tree_add_106_2_groupi_n_941) | (csa_tree_add_106_2_groupi_n_941
    & csa_tree_add_106_2_groupi_n_987)));
 assign csa_tree_add_106_2_groupi_n_1052 = (csa_tree_add_106_2_groupi_n_1015 ^ (csa_tree_add_106_2_groupi_n_941
    ^ csa_tree_add_106_2_groupi_n_987));
 assign csa_tree_add_106_2_groupi_n_1049 = ((csa_tree_add_106_2_groupi_n_1001 & csa_tree_add_106_2_groupi_n_839)
    | ((csa_tree_add_106_2_groupi_n_839 & csa_tree_add_106_2_groupi_n_907) | (csa_tree_add_106_2_groupi_n_907
    & csa_tree_add_106_2_groupi_n_1001)));
 assign csa_tree_add_106_2_groupi_n_1050 = (csa_tree_add_106_2_groupi_n_839 ^ (csa_tree_add_106_2_groupi_n_907
    ^ csa_tree_add_106_2_groupi_n_1001));
 assign csa_tree_add_106_2_groupi_n_1047 = ((csa_tree_add_106_2_groupi_n_999 & csa_tree_add_106_2_groupi_n_364)
    | ((csa_tree_add_106_2_groupi_n_364 & csa_tree_add_106_2_groupi_n_452) | (csa_tree_add_106_2_groupi_n_452
    & csa_tree_add_106_2_groupi_n_999)));
 assign csa_tree_add_106_2_groupi_n_1048 = (csa_tree_add_106_2_groupi_n_364 ^ (csa_tree_add_106_2_groupi_n_452
    ^ csa_tree_add_106_2_groupi_n_999));
 assign csa_tree_add_106_2_groupi_n_1043 = ((csa_tree_add_106_2_groupi_n_985 & csa_tree_add_106_2_groupi_n_449)
    | ((csa_tree_add_106_2_groupi_n_449 & csa_tree_add_106_2_groupi_n_980) | (csa_tree_add_106_2_groupi_n_980
    & csa_tree_add_106_2_groupi_n_985)));
 assign csa_tree_add_106_2_groupi_n_1044 = (csa_tree_add_106_2_groupi_n_449 ^ (csa_tree_add_106_2_groupi_n_980
    ^ csa_tree_add_106_2_groupi_n_985));
 assign csa_tree_add_106_2_groupi_n_1041 = ((csa_tree_add_106_2_groupi_n_1000 & csa_tree_add_106_2_groupi_n_970)
    | ((csa_tree_add_106_2_groupi_n_970 & csa_tree_add_106_2_groupi_n_877) | (csa_tree_add_106_2_groupi_n_877
    & csa_tree_add_106_2_groupi_n_1000)));
 assign csa_tree_add_106_2_groupi_n_1042 = (csa_tree_add_106_2_groupi_n_970 ^ (csa_tree_add_106_2_groupi_n_877
    ^ csa_tree_add_106_2_groupi_n_1000));
 assign csa_tree_add_106_2_groupi_n_1039 = ((csa_tree_add_106_2_groupi_n_1009 & csa_tree_add_106_2_groupi_n_381)
    | ((csa_tree_add_106_2_groupi_n_381 & csa_tree_add_106_2_groupi_n_971) | (csa_tree_add_106_2_groupi_n_971
    & csa_tree_add_106_2_groupi_n_1009)));
 assign csa_tree_add_106_2_groupi_n_1040 = (csa_tree_add_106_2_groupi_n_381 ^ (csa_tree_add_106_2_groupi_n_971
    ^ csa_tree_add_106_2_groupi_n_1009));
 assign csa_tree_add_106_2_groupi_n_1038 = ~(csa_tree_add_106_2_groupi_n_1013 ^ csa_tree_add_106_2_groupi_n_1003);
 assign csa_tree_add_106_2_groupi_n_1034 = ((csa_tree_add_106_2_groupi_n_935 & csa_tree_add_106_2_groupi_n_876)
    | ((csa_tree_add_106_2_groupi_n_876 & csa_tree_add_106_2_groupi_n_959) | (csa_tree_add_106_2_groupi_n_959
    & csa_tree_add_106_2_groupi_n_935)));
 assign csa_tree_add_106_2_groupi_n_1035 = (csa_tree_add_106_2_groupi_n_876 ^ (csa_tree_add_106_2_groupi_n_959
    ^ csa_tree_add_106_2_groupi_n_935));
 assign csa_tree_add_106_2_groupi_n_1030 = ((csa_tree_add_106_2_groupi_n_984 & csa_tree_add_106_2_groupi_n_521)
    | ((csa_tree_add_106_2_groupi_n_521 & csa_tree_add_106_2_groupi_n_792) | (csa_tree_add_106_2_groupi_n_792
    & csa_tree_add_106_2_groupi_n_984)));
 assign csa_tree_add_106_2_groupi_n_1031 = (csa_tree_add_106_2_groupi_n_521 ^ (csa_tree_add_106_2_groupi_n_792
    ^ csa_tree_add_106_2_groupi_n_984));
 assign csa_tree_add_106_2_groupi_n_1028 = ((csa_tree_add_106_2_groupi_n_960 & csa_tree_add_106_2_groupi_n_512)
    | ((csa_tree_add_106_2_groupi_n_512 & csa_tree_add_106_2_groupi_n_903) | (csa_tree_add_106_2_groupi_n_903
    & csa_tree_add_106_2_groupi_n_960)));
 assign csa_tree_add_106_2_groupi_n_1029 = (csa_tree_add_106_2_groupi_n_512 ^ (csa_tree_add_106_2_groupi_n_903
    ^ csa_tree_add_106_2_groupi_n_960));
 assign csa_tree_add_106_2_groupi_n_1024 = ((csa_tree_add_106_2_groupi_n_958 & csa_tree_add_106_2_groupi_n_506)
    | ((csa_tree_add_106_2_groupi_n_506 & csa_tree_add_106_2_groupi_n_746) | (csa_tree_add_106_2_groupi_n_746
    & csa_tree_add_106_2_groupi_n_958)));
 assign csa_tree_add_106_2_groupi_n_1025 = (csa_tree_add_106_2_groupi_n_506 ^ (csa_tree_add_106_2_groupi_n_746
    ^ csa_tree_add_106_2_groupi_n_958));
 assign csa_tree_add_106_2_groupi_n_1022 = ((csa_tree_add_106_2_groupi_n_982 & csa_tree_add_106_2_groupi_n_693)
    | ((csa_tree_add_106_2_groupi_n_693 & csa_tree_add_106_2_groupi_n_936) | (csa_tree_add_106_2_groupi_n_936
    & csa_tree_add_106_2_groupi_n_982)));
 assign csa_tree_add_106_2_groupi_n_1023 = (csa_tree_add_106_2_groupi_n_693 ^ (csa_tree_add_106_2_groupi_n_936
    ^ csa_tree_add_106_2_groupi_n_982));
 assign csa_tree_add_106_2_groupi_n_1020 = ((csa_tree_add_106_2_groupi_n_961 & csa_tree_add_106_2_groupi_n_436)
    | ((csa_tree_add_106_2_groupi_n_436 & csa_tree_add_106_2_groupi_n_934) | (csa_tree_add_106_2_groupi_n_934
    & csa_tree_add_106_2_groupi_n_961)));
 assign csa_tree_add_106_2_groupi_n_1021 = (csa_tree_add_106_2_groupi_n_436 ^ (csa_tree_add_106_2_groupi_n_934
    ^ csa_tree_add_106_2_groupi_n_961));
 assign csa_tree_add_106_2_groupi_n_1018 = ((csa_tree_add_106_2_groupi_n_956 & csa_tree_add_106_2_groupi_n_925)
    | ((csa_tree_add_106_2_groupi_n_925 & csa_tree_add_106_2_groupi_n_905) | (csa_tree_add_106_2_groupi_n_905
    & csa_tree_add_106_2_groupi_n_956)));
 assign csa_tree_add_106_2_groupi_n_1019 = (csa_tree_add_106_2_groupi_n_925 ^ (csa_tree_add_106_2_groupi_n_905
    ^ csa_tree_add_106_2_groupi_n_956));
 assign csa_tree_add_106_2_groupi_n_1014 = ((csa_tree_add_106_2_groupi_n_917 & csa_tree_add_106_2_groupi_n_382)
    | ((csa_tree_add_106_2_groupi_n_382 & csa_tree_add_106_2_groupi_n_964) | (csa_tree_add_106_2_groupi_n_964
    & csa_tree_add_106_2_groupi_n_917)));
 assign csa_tree_add_106_2_groupi_n_1015 = (csa_tree_add_106_2_groupi_n_382 ^ (csa_tree_add_106_2_groupi_n_964
    ^ csa_tree_add_106_2_groupi_n_917));
 assign csa_tree_add_106_2_groupi_n_1013 = ~(csa_tree_add_106_2_groupi_n_986 ^ csa_tree_add_106_2_groupi_n_927);
 assign csa_tree_add_106_2_groupi_n_1009 = ((csa_tree_add_106_2_groupi_n_969 & csa_tree_add_106_2_groupi_n_380)
    | ((csa_tree_add_106_2_groupi_n_380 & csa_tree_add_106_2_groupi_n_931) | (csa_tree_add_106_2_groupi_n_931
    & csa_tree_add_106_2_groupi_n_969)));
 assign csa_tree_add_106_2_groupi_n_1010 = (csa_tree_add_106_2_groupi_n_380 ^ (csa_tree_add_106_2_groupi_n_931
    ^ csa_tree_add_106_2_groupi_n_969));
 assign csa_tree_add_106_2_groupi_n_1007 = ((csa_tree_add_106_2_groupi_n_968 & csa_tree_add_106_2_groupi_n_450)
    | ((csa_tree_add_106_2_groupi_n_450 & csa_tree_add_106_2_groupi_n_933) | (csa_tree_add_106_2_groupi_n_933
    & csa_tree_add_106_2_groupi_n_968)));
 assign csa_tree_add_106_2_groupi_n_1008 = (csa_tree_add_106_2_groupi_n_450 ^ (csa_tree_add_106_2_groupi_n_933
    ^ csa_tree_add_106_2_groupi_n_968));
 assign csa_tree_add_106_2_groupi_n_1005 = ((csa_tree_add_106_2_groupi_n_966 & csa_tree_add_106_2_groupi_n_914)
    | ((csa_tree_add_106_2_groupi_n_914 & csa_tree_add_106_2_groupi_n_899) | (csa_tree_add_106_2_groupi_n_899
    & csa_tree_add_106_2_groupi_n_966)));
 assign csa_tree_add_106_2_groupi_n_1006 = (csa_tree_add_106_2_groupi_n_914 ^ (csa_tree_add_106_2_groupi_n_899
    ^ csa_tree_add_106_2_groupi_n_966));
 assign csa_tree_add_106_2_groupi_n_1003 = ((csa_tree_add_106_2_groupi_n_962 & csa_tree_add_106_2_groupi_n_870)
    | ((csa_tree_add_106_2_groupi_n_870 & csa_tree_add_106_2_groupi_n_881) | (csa_tree_add_106_2_groupi_n_881
    & csa_tree_add_106_2_groupi_n_962)));
 assign csa_tree_add_106_2_groupi_n_1004 = (csa_tree_add_106_2_groupi_n_870 ^ (csa_tree_add_106_2_groupi_n_881
    ^ csa_tree_add_106_2_groupi_n_962));
 assign csa_tree_add_106_2_groupi_n_1001 = ((csa_tree_add_106_2_groupi_n_938 & csa_tree_add_106_2_groupi_n_375)
    | ((csa_tree_add_106_2_groupi_n_375 & csa_tree_add_106_2_groupi_n_435) | (csa_tree_add_106_2_groupi_n_435
    & csa_tree_add_106_2_groupi_n_938)));
 assign csa_tree_add_106_2_groupi_n_1002 = (csa_tree_add_106_2_groupi_n_375 ^ (csa_tree_add_106_2_groupi_n_435
    ^ csa_tree_add_106_2_groupi_n_938));
 assign csa_tree_add_106_2_groupi_n_999 = ((csa_tree_add_106_2_groupi_n_932 & csa_tree_add_106_2_groupi_n_442)
    | ((csa_tree_add_106_2_groupi_n_442 & csa_tree_add_106_2_groupi_n_921) | (csa_tree_add_106_2_groupi_n_921
    & csa_tree_add_106_2_groupi_n_932)));
 assign csa_tree_add_106_2_groupi_n_1000 = (csa_tree_add_106_2_groupi_n_442 ^ (csa_tree_add_106_2_groupi_n_921
    ^ csa_tree_add_106_2_groupi_n_932));
 assign csa_tree_add_106_2_groupi_n_993 = ((csa_tree_add_106_2_groupi_n_915 & csa_tree_add_106_2_groupi_n_383)
    | ((csa_tree_add_106_2_groupi_n_383 & csa_tree_add_106_2_groupi_n_942) | (csa_tree_add_106_2_groupi_n_942
    & csa_tree_add_106_2_groupi_n_915)));
 assign csa_tree_add_106_2_groupi_n_994 = (csa_tree_add_106_2_groupi_n_383 ^ (csa_tree_add_106_2_groupi_n_942
    ^ csa_tree_add_106_2_groupi_n_915));
 assign csa_tree_add_106_2_groupi_n_991 = ((csa_tree_add_106_2_groupi_n_895 & csa_tree_add_106_2_groupi_n_916)
    | ((csa_tree_add_106_2_groupi_n_916 & csa_tree_add_106_2_groupi_n_940) | (csa_tree_add_106_2_groupi_n_940
    & csa_tree_add_106_2_groupi_n_895)));
 assign csa_tree_add_106_2_groupi_n_992 = (csa_tree_add_106_2_groupi_n_916 ^ (csa_tree_add_106_2_groupi_n_940
    ^ csa_tree_add_106_2_groupi_n_895));
 assign csa_tree_add_106_2_groupi_n_987 = ((csa_tree_add_106_2_groupi_n_946 & csa_tree_add_106_2_groupi_n_376)
    | ((csa_tree_add_106_2_groupi_n_376 & csa_tree_add_106_2_groupi_n_893) | (csa_tree_add_106_2_groupi_n_893
    & csa_tree_add_106_2_groupi_n_946)));
 assign csa_tree_add_106_2_groupi_n_988 = (csa_tree_add_106_2_groupi_n_376 ^ (csa_tree_add_106_2_groupi_n_893
    ^ csa_tree_add_106_2_groupi_n_946));
 assign csa_tree_add_106_2_groupi_n_986 = ~(csa_tree_add_106_2_groupi_n_926 ^ csa_tree_add_106_2_groupi_n_972);
 assign csa_tree_add_106_2_groupi_n_984 = ((csa_tree_add_106_2_groupi_n_944 & csa_tree_add_106_2_groupi_n_567)
    | ((csa_tree_add_106_2_groupi_n_567 & csa_tree_add_106_2_groupi_n_758) | (csa_tree_add_106_2_groupi_n_758
    & csa_tree_add_106_2_groupi_n_944)));
 assign csa_tree_add_106_2_groupi_n_985 = (csa_tree_add_106_2_groupi_n_567 ^ (csa_tree_add_106_2_groupi_n_758
    ^ csa_tree_add_106_2_groupi_n_944));
 assign csa_tree_add_106_2_groupi_n_980 = ((csa_tree_add_106_2_groupi_n_945 & csa_tree_add_106_2_groupi_n_499)
    | ((csa_tree_add_106_2_groupi_n_499 & csa_tree_add_106_2_groupi_n_832) | (csa_tree_add_106_2_groupi_n_832
    & csa_tree_add_106_2_groupi_n_945)));
 assign csa_tree_add_106_2_groupi_n_981 = (csa_tree_add_106_2_groupi_n_499 ^ (csa_tree_add_106_2_groupi_n_832
    ^ csa_tree_add_106_2_groupi_n_945));
 assign csa_tree_add_106_2_groupi_n_976 = ((csa_tree_add_106_2_groupi_n_904 & csa_tree_add_106_2_groupi_n_374)
    | ((csa_tree_add_106_2_groupi_n_374 & csa_tree_add_106_2_groupi_n_873) | (csa_tree_add_106_2_groupi_n_873
    & csa_tree_add_106_2_groupi_n_904)));
 assign csa_tree_add_106_2_groupi_n_977 = (csa_tree_add_106_2_groupi_n_374 ^ (csa_tree_add_106_2_groupi_n_873
    ^ csa_tree_add_106_2_groupi_n_904));
 assign csa_tree_add_106_2_groupi_n_974 = ((csa_tree_add_106_2_groupi_n_898 & csa_tree_add_106_2_groupi_n_372)
    | ((csa_tree_add_106_2_groupi_n_372 & csa_tree_add_106_2_groupi_n_884) | (csa_tree_add_106_2_groupi_n_884
    & csa_tree_add_106_2_groupi_n_898)));
 assign csa_tree_add_106_2_groupi_n_975 = (csa_tree_add_106_2_groupi_n_372 ^ (csa_tree_add_106_2_groupi_n_884
    ^ csa_tree_add_106_2_groupi_n_898));
 assign csa_tree_add_106_2_groupi_n_966 = ((csa_tree_add_106_2_groupi_n_894 & csa_tree_add_106_2_groupi_n_879)
    | ((csa_tree_add_106_2_groupi_n_879 & csa_tree_add_106_2_groupi_n_874) | (csa_tree_add_106_2_groupi_n_874
    & csa_tree_add_106_2_groupi_n_894)));
 assign csa_tree_add_106_2_groupi_n_967 = (csa_tree_add_106_2_groupi_n_879 ^ (csa_tree_add_106_2_groupi_n_874
    ^ csa_tree_add_106_2_groupi_n_894));
 assign csa_tree_add_106_2_groupi_n_964 = ((csa_tree_add_106_2_groupi_n_928 & csa_tree_add_106_2_groupi_n_843)
    | ((csa_tree_add_106_2_groupi_n_843 & csa_tree_add_106_2_groupi_n_840) | (csa_tree_add_106_2_groupi_n_840
    & csa_tree_add_106_2_groupi_n_928)));
 assign csa_tree_add_106_2_groupi_n_965 = (csa_tree_add_106_2_groupi_n_843 ^ (csa_tree_add_106_2_groupi_n_840
    ^ csa_tree_add_106_2_groupi_n_928));
 assign csa_tree_add_106_2_groupi_n_960 = ((csa_tree_add_106_2_groupi_n_882 & csa_tree_add_106_2_groupi_n_574)
    | ((csa_tree_add_106_2_groupi_n_574 & csa_tree_add_106_2_groupi_n_853) | (csa_tree_add_106_2_groupi_n_853
    & csa_tree_add_106_2_groupi_n_882)));
 assign csa_tree_add_106_2_groupi_n_961 = (csa_tree_add_106_2_groupi_n_574 ^ (csa_tree_add_106_2_groupi_n_853
    ^ csa_tree_add_106_2_groupi_n_882));
 assign csa_tree_add_106_2_groupi_n_956 = ((csa_tree_add_106_2_groupi_n_878 & csa_tree_add_106_2_groupi_n_365)
    | ((csa_tree_add_106_2_groupi_n_365 & csa_tree_add_106_2_groupi_n_885) | (csa_tree_add_106_2_groupi_n_885
    & csa_tree_add_106_2_groupi_n_878)));
 assign csa_tree_add_106_2_groupi_n_957 = (csa_tree_add_106_2_groupi_n_365 ^ (csa_tree_add_106_2_groupi_n_885
    ^ csa_tree_add_106_2_groupi_n_878));
 assign csa_tree_add_106_2_groupi_n_946 = ((csa_tree_add_106_2_groupi_n_906 & csa_tree_add_106_2_groupi_n_841)
    | ((csa_tree_add_106_2_groupi_n_841 & csa_tree_add_106_2_groupi_n_796) | (csa_tree_add_106_2_groupi_n_796
    & csa_tree_add_106_2_groupi_n_906)));
 assign csa_tree_add_106_2_groupi_n_947 = (csa_tree_add_106_2_groupi_n_841 ^ (csa_tree_add_106_2_groupi_n_796
    ^ csa_tree_add_106_2_groupi_n_906));
 assign csa_tree_add_106_2_groupi_n_944 = ((csa_tree_add_106_2_groupi_n_902 & csa_tree_add_106_2_groupi_n_566)
    | ((csa_tree_add_106_2_groupi_n_566 & csa_tree_add_106_2_groupi_n_679) | (csa_tree_add_106_2_groupi_n_679
    & csa_tree_add_106_2_groupi_n_902)));
 assign csa_tree_add_106_2_groupi_n_945 = (csa_tree_add_106_2_groupi_n_566 ^ (csa_tree_add_106_2_groupi_n_679
    ^ csa_tree_add_106_2_groupi_n_902));
 assign csa_tree_add_106_2_groupi_n_942 = ((csa_tree_add_106_2_groupi_n_875 & csa_tree_add_106_2_groupi_n_373)
    | ((csa_tree_add_106_2_groupi_n_373 & csa_tree_add_106_2_groupi_n_844) | (csa_tree_add_106_2_groupi_n_844
    & csa_tree_add_106_2_groupi_n_875)));
 assign csa_tree_add_106_2_groupi_n_943 = (csa_tree_add_106_2_groupi_n_373 ^ (csa_tree_add_106_2_groupi_n_844
    ^ csa_tree_add_106_2_groupi_n_875));
 assign csa_tree_add_106_2_groupi_n_940 = ((csa_tree_add_106_2_groupi_n_892 & csa_tree_add_106_2_groupi_n_457)
    | ((csa_tree_add_106_2_groupi_n_457 & csa_tree_add_106_2_groupi_n_845) | (csa_tree_add_106_2_groupi_n_845
    & csa_tree_add_106_2_groupi_n_892)));
 assign csa_tree_add_106_2_groupi_n_941 = (csa_tree_add_106_2_groupi_n_457 ^ (csa_tree_add_106_2_groupi_n_845
    ^ csa_tree_add_106_2_groupi_n_892));
 assign csa_tree_add_106_2_groupi_n_938 = ((csa_tree_add_106_2_groupi_n_850 & csa_tree_add_106_2_groupi_n_515)
    | ((csa_tree_add_106_2_groupi_n_515 & csa_tree_add_106_2_groupi_n_802) | (csa_tree_add_106_2_groupi_n_802
    & csa_tree_add_106_2_groupi_n_850)));
 assign csa_tree_add_106_2_groupi_n_939 = (csa_tree_add_106_2_groupi_n_515 ^ (csa_tree_add_106_2_groupi_n_802
    ^ csa_tree_add_106_2_groupi_n_850));
 assign csa_tree_add_106_2_groupi_n_934 = ((csa_tree_add_106_2_groupi_n_883 & csa_tree_add_106_2_groupi_n_556)
    | ((csa_tree_add_106_2_groupi_n_556 & csa_tree_add_106_2_groupi_n_500) | (csa_tree_add_106_2_groupi_n_500
    & csa_tree_add_106_2_groupi_n_883)));
 assign csa_tree_add_106_2_groupi_n_935 = (csa_tree_add_106_2_groupi_n_556 ^ (csa_tree_add_106_2_groupi_n_500
    ^ csa_tree_add_106_2_groupi_n_883));
 assign csa_tree_add_106_2_groupi_n_928 = ((csa_tree_add_106_2_groupi_n_838 & csa_tree_add_106_2_groupi_n_458)
    | ((csa_tree_add_106_2_groupi_n_458 & csa_tree_add_106_2_groupi_n_527) | (csa_tree_add_106_2_groupi_n_527
    & csa_tree_add_106_2_groupi_n_838)));
 assign csa_tree_add_106_2_groupi_n_929 = (csa_tree_add_106_2_groupi_n_458 ^ (csa_tree_add_106_2_groupi_n_527
    ^ csa_tree_add_106_2_groupi_n_838));
 assign csa_tree_add_106_2_groupi_n_927 = ~(csa_tree_add_106_2_groupi_n_886 ^ csa_tree_add_106_2_groupi_n_880);
 assign csa_tree_add_106_2_groupi_n_924 = ((csa_tree_add_106_2_groupi_n_823 & csa_tree_add_106_2_groupi_n_448)
    | ((csa_tree_add_106_2_groupi_n_448 & csa_tree_add_106_2_groupi_n_507) | (csa_tree_add_106_2_groupi_n_507
    & csa_tree_add_106_2_groupi_n_823)));
 assign csa_tree_add_106_2_groupi_n_925 = (csa_tree_add_106_2_groupi_n_448 ^ (csa_tree_add_106_2_groupi_n_507
    ^ csa_tree_add_106_2_groupi_n_823));
 assign csa_tree_add_106_2_groupi_n_916 = ((csa_tree_add_106_2_groupi_n_842 & csa_tree_add_106_2_groupi_n_811)
    | ((csa_tree_add_106_2_groupi_n_811 & csa_tree_add_106_2_groupi_n_816) | (csa_tree_add_106_2_groupi_n_816
    & csa_tree_add_106_2_groupi_n_842)));
 assign csa_tree_add_106_2_groupi_n_917 = (csa_tree_add_106_2_groupi_n_811 ^ (csa_tree_add_106_2_groupi_n_816
    ^ csa_tree_add_106_2_groupi_n_842));
 assign csa_tree_add_106_2_groupi_n_914 = ((csa_tree_add_106_2_groupi_n_835 & csa_tree_add_106_2_groupi_n_441)
    | ((csa_tree_add_106_2_groupi_n_441 & csa_tree_add_106_2_groupi_n_488) | (csa_tree_add_106_2_groupi_n_488
    & csa_tree_add_106_2_groupi_n_835)));
 assign csa_tree_add_106_2_groupi_n_915 = (csa_tree_add_106_2_groupi_n_441 ^ (csa_tree_add_106_2_groupi_n_488
    ^ csa_tree_add_106_2_groupi_n_835));
 assign csa_tree_add_106_2_groupi_n_906 = ((csa_tree_add_106_2_groupi_n_856 & csa_tree_add_106_2_groupi_n_524)
    | ((csa_tree_add_106_2_groupi_n_524 & csa_tree_add_106_2_groupi_n_785) | (csa_tree_add_106_2_groupi_n_785
    & csa_tree_add_106_2_groupi_n_856)));
 assign csa_tree_add_106_2_groupi_n_907 = (csa_tree_add_106_2_groupi_n_524 ^ (csa_tree_add_106_2_groupi_n_785
    ^ csa_tree_add_106_2_groupi_n_856));
 assign csa_tree_add_106_2_groupi_n_904 = ((csa_tree_add_106_2_groupi_n_819 & csa_tree_add_106_2_groupi_n_559)
    | ((csa_tree_add_106_2_groupi_n_559 & csa_tree_add_106_2_groupi_n_781) | (csa_tree_add_106_2_groupi_n_781
    & csa_tree_add_106_2_groupi_n_819)));
 assign csa_tree_add_106_2_groupi_n_905 = (csa_tree_add_106_2_groupi_n_559 ^ (csa_tree_add_106_2_groupi_n_781
    ^ csa_tree_add_106_2_groupi_n_819));
 assign csa_tree_add_106_2_groupi_n_902 = ((csa_tree_add_106_2_groupi_n_852 & csa_tree_add_106_2_groupi_n_477)
    | ((csa_tree_add_106_2_groupi_n_477 & csa_tree_add_106_2_groupi_n_565) | (csa_tree_add_106_2_groupi_n_565
    & csa_tree_add_106_2_groupi_n_852)));
 assign csa_tree_add_106_2_groupi_n_903 = (csa_tree_add_106_2_groupi_n_477 ^ (csa_tree_add_106_2_groupi_n_565
    ^ csa_tree_add_106_2_groupi_n_852));
 assign csa_tree_add_106_2_groupi_n_898 = ((csa_tree_add_106_2_groupi_n_820 & csa_tree_add_106_2_groupi_n_443)
    | ((csa_tree_add_106_2_groupi_n_443 & csa_tree_add_106_2_groupi_n_490) | (csa_tree_add_106_2_groupi_n_490
    & csa_tree_add_106_2_groupi_n_820)));
 assign csa_tree_add_106_2_groupi_n_899 = (csa_tree_add_106_2_groupi_n_443 ^ (csa_tree_add_106_2_groupi_n_490
    ^ csa_tree_add_106_2_groupi_n_820));
 assign csa_tree_add_106_2_groupi_n_894 = ((csa_tree_add_106_2_groupi_n_814 & csa_tree_add_106_2_groupi_n_447)
    | ((csa_tree_add_106_2_groupi_n_447 & csa_tree_add_106_2_groupi_n_492) | (csa_tree_add_106_2_groupi_n_492
    & csa_tree_add_106_2_groupi_n_814)));
 assign csa_tree_add_106_2_groupi_n_895 = (csa_tree_add_106_2_groupi_n_447 ^ (csa_tree_add_106_2_groupi_n_492
    ^ csa_tree_add_106_2_groupi_n_814));
 assign csa_tree_add_106_2_groupi_n_892 = ((csa_tree_add_106_2_groupi_n_812 & csa_tree_add_106_2_groupi_n_440)
    | ((csa_tree_add_106_2_groupi_n_440 & csa_tree_add_106_2_groupi_n_502) | (csa_tree_add_106_2_groupi_n_502
    & csa_tree_add_106_2_groupi_n_812)));
 assign csa_tree_add_106_2_groupi_n_893 = (csa_tree_add_106_2_groupi_n_440 ^ (csa_tree_add_106_2_groupi_n_502
    ^ csa_tree_add_106_2_groupi_n_812));
 assign csa_tree_add_106_2_groupi_n_888 = ((csa_tree_add_106_2_groupi_n_808 & csa_tree_add_106_2_groupi_n_453)
    | ((csa_tree_add_106_2_groupi_n_453 & csa_tree_add_106_2_groupi_n_517) | (csa_tree_add_106_2_groupi_n_517
    & csa_tree_add_106_2_groupi_n_808)));
 assign csa_tree_add_106_2_groupi_n_889 = (csa_tree_add_106_2_groupi_n_453 ^ (csa_tree_add_106_2_groupi_n_517
    ^ csa_tree_add_106_2_groupi_n_808));
 assign csa_tree_add_106_2_groupi_n_884 = ((csa_tree_add_106_2_groupi_n_834 & csa_tree_add_106_2_groupi_n_543)
    | ((csa_tree_add_106_2_groupi_n_543 & csa_tree_add_106_2_groupi_n_789) | (csa_tree_add_106_2_groupi_n_789
    & csa_tree_add_106_2_groupi_n_834)));
 assign csa_tree_add_106_2_groupi_n_885 = (csa_tree_add_106_2_groupi_n_543 ^ (csa_tree_add_106_2_groupi_n_789
    ^ csa_tree_add_106_2_groupi_n_834));
 assign csa_tree_add_106_2_groupi_n_882 = ((csa_tree_add_106_2_groupi_n_797 & csa_tree_add_106_2_groupi_n_555)
    | ((csa_tree_add_106_2_groupi_n_555 & csa_tree_add_106_2_groupi_n_510) | (csa_tree_add_106_2_groupi_n_510
    & csa_tree_add_106_2_groupi_n_797)));
 assign csa_tree_add_106_2_groupi_n_883 = (csa_tree_add_106_2_groupi_n_555 ^ (csa_tree_add_106_2_groupi_n_510
    ^ csa_tree_add_106_2_groupi_n_797));
 assign csa_tree_add_106_2_groupi_n_878 = ((csa_tree_add_106_2_groupi_n_813 & csa_tree_add_106_2_groupi_n_546)
    | ((csa_tree_add_106_2_groupi_n_546 & csa_tree_add_106_2_groupi_n_786) | (csa_tree_add_106_2_groupi_n_786
    & csa_tree_add_106_2_groupi_n_813)));
 assign csa_tree_add_106_2_groupi_n_879 = (csa_tree_add_106_2_groupi_n_546 ^ (csa_tree_add_106_2_groupi_n_786
    ^ csa_tree_add_106_2_groupi_n_813));
 assign csa_tree_add_106_2_groupi_n_876 = ((csa_tree_add_106_2_groupi_n_798 & csa_tree_add_106_2_groupi_n_590)
    | ((csa_tree_add_106_2_groupi_n_590 & csa_tree_add_106_2_groupi_n_489) | (csa_tree_add_106_2_groupi_n_489
    & csa_tree_add_106_2_groupi_n_798)));
 assign csa_tree_add_106_2_groupi_n_877 = (csa_tree_add_106_2_groupi_n_590 ^ (csa_tree_add_106_2_groupi_n_489
    ^ csa_tree_add_106_2_groupi_n_798));
 assign csa_tree_add_106_2_groupi_n_874 = ((csa_tree_add_106_2_groupi_n_815 & csa_tree_add_106_2_groupi_n_562)
    | ((csa_tree_add_106_2_groupi_n_562 & csa_tree_add_106_2_groupi_n_787) | (csa_tree_add_106_2_groupi_n_787
    & csa_tree_add_106_2_groupi_n_815)));
 assign csa_tree_add_106_2_groupi_n_875 = (csa_tree_add_106_2_groupi_n_562 ^ (csa_tree_add_106_2_groupi_n_787
    ^ csa_tree_add_106_2_groupi_n_815));
 assign csa_tree_add_106_2_groupi_n_872 = ((csa_tree_add_106_2_groupi_n_822 & csa_tree_add_106_2_groupi_n_569)
    | ((csa_tree_add_106_2_groupi_n_569 & csa_tree_add_106_2_groupi_n_744) | (csa_tree_add_106_2_groupi_n_744
    & csa_tree_add_106_2_groupi_n_822)));
 assign csa_tree_add_106_2_groupi_n_873 = (csa_tree_add_106_2_groupi_n_569 ^ (csa_tree_add_106_2_groupi_n_744
    ^ csa_tree_add_106_2_groupi_n_822));
 assign csa_tree_add_106_2_groupi_n_856 = ((csa_tree_add_106_2_groupi_n_801 & csa_tree_add_106_2_groupi_n_573)
    | ((csa_tree_add_106_2_groupi_n_573 & csa_tree_add_106_2_groupi_n_734) | (csa_tree_add_106_2_groupi_n_734
    & csa_tree_add_106_2_groupi_n_801)));
 assign csa_tree_add_106_2_groupi_n_857 = (csa_tree_add_106_2_groupi_n_573 ^ (csa_tree_add_106_2_groupi_n_734
    ^ csa_tree_add_106_2_groupi_n_801));
 assign csa_tree_add_106_2_groupi_n_855 = ~(csa_tree_add_106_2_groupi_n_427 ^ csa_tree_add_106_2_groupi_n_830);
 assign csa_tree_add_106_2_groupi_n_854 = ~(csa_tree_add_106_2_groupi_n_0 ^ csa_tree_add_106_2_groupi_n_821);
 assign csa_tree_add_106_2_groupi_n_850 = ((csa_tree_add_106_2_groupi_n_769 & csa_tree_add_106_2_groupi_n_568)
    | ((csa_tree_add_106_2_groupi_n_568 & csa_tree_add_106_2_groupi_n_763) | (csa_tree_add_106_2_groupi_n_763
    & csa_tree_add_106_2_groupi_n_769)));
 assign csa_tree_add_106_2_groupi_n_851 = (csa_tree_add_106_2_groupi_n_568 ^ (csa_tree_add_106_2_groupi_n_763
    ^ csa_tree_add_106_2_groupi_n_769));
 assign csa_tree_add_106_2_groupi_n_844 = ((csa_tree_add_106_2_groupi_n_773 & csa_tree_add_106_2_groupi_n_484)
    | ((csa_tree_add_106_2_groupi_n_484 & csa_tree_add_106_2_groupi_n_550) | (csa_tree_add_106_2_groupi_n_550
    & csa_tree_add_106_2_groupi_n_773)));
 assign csa_tree_add_106_2_groupi_n_845 = (csa_tree_add_106_2_groupi_n_484 ^ (csa_tree_add_106_2_groupi_n_550
    ^ csa_tree_add_106_2_groupi_n_773));
 assign csa_tree_add_106_2_groupi_n_842 = ((csa_tree_add_106_2_groupi_n_795 & csa_tree_add_106_2_groupi_n_549)
    | ((csa_tree_add_106_2_groupi_n_549 & csa_tree_add_106_2_groupi_n_685) | (csa_tree_add_106_2_groupi_n_685
    & csa_tree_add_106_2_groupi_n_795)));
 assign csa_tree_add_106_2_groupi_n_843 = (csa_tree_add_106_2_groupi_n_549 ^ (csa_tree_add_106_2_groupi_n_685
    ^ csa_tree_add_106_2_groupi_n_795));
 assign csa_tree_add_106_2_groupi_n_840 = ((csa_tree_add_106_2_groupi_n_775 & csa_tree_add_106_2_groupi_n_583)
    | ((csa_tree_add_106_2_groupi_n_583 & csa_tree_add_106_2_groupi_n_784) | (csa_tree_add_106_2_groupi_n_784
    & csa_tree_add_106_2_groupi_n_775)));
 assign csa_tree_add_106_2_groupi_n_841 = (csa_tree_add_106_2_groupi_n_583 ^ (csa_tree_add_106_2_groupi_n_784
    ^ csa_tree_add_106_2_groupi_n_775));
 assign csa_tree_add_106_2_groupi_n_838 = ((csa_tree_add_106_2_groupi_n_791 & csa_tree_add_106_2_groupi_n_578)
    | ((csa_tree_add_106_2_groupi_n_578 & csa_tree_add_106_2_groupi_n_724) | (csa_tree_add_106_2_groupi_n_724
    & csa_tree_add_106_2_groupi_n_791)));
 assign csa_tree_add_106_2_groupi_n_839 = (csa_tree_add_106_2_groupi_n_578 ^ (csa_tree_add_106_2_groupi_n_724
    ^ csa_tree_add_106_2_groupi_n_791));
 assign csa_tree_add_106_2_groupi_n_834 = ((csa_tree_add_106_2_groupi_n_783 & csa_tree_add_106_2_groupi_n_394)
    | ((csa_tree_add_106_2_groupi_n_394 & csa_tree_add_106_2_groupi_n_754) | (csa_tree_add_106_2_groupi_n_754
    & csa_tree_add_106_2_groupi_n_783)));
 assign csa_tree_add_106_2_groupi_n_835 = (csa_tree_add_106_2_groupi_n_394 ^ (csa_tree_add_106_2_groupi_n_754
    ^ csa_tree_add_106_2_groupi_n_783));
 assign csa_tree_add_106_2_groupi_n_832 = ((csa_tree_add_106_2_groupi_n_764 & csa_tree_add_106_2_groupi_n_588)
    | ((csa_tree_add_106_2_groupi_n_588 & csa_tree_add_106_2_groupi_n_745) | (csa_tree_add_106_2_groupi_n_745
    & csa_tree_add_106_2_groupi_n_764)));
 assign csa_tree_add_106_2_groupi_n_833 = (csa_tree_add_106_2_groupi_n_588 ^ (csa_tree_add_106_2_groupi_n_745
    ^ csa_tree_add_106_2_groupi_n_764));
 assign csa_tree_add_106_2_groupi_n_824 = ((csa_tree_add_106_2_groupi_n_737 & csa_tree_add_106_2_groupi_n_777)
    | ((csa_tree_add_106_2_groupi_n_777 & csa_tree_add_106_2_groupi_n_701) | (csa_tree_add_106_2_groupi_n_701
    & csa_tree_add_106_2_groupi_n_737)));
 assign csa_tree_add_106_2_groupi_n_825 = (csa_tree_add_106_2_groupi_n_777 ^ (csa_tree_add_106_2_groupi_n_701
    ^ csa_tree_add_106_2_groupi_n_737));
 assign csa_tree_add_106_2_groupi_n_822 = ((csa_tree_add_106_2_groupi_n_788 & csa_tree_add_106_2_groupi_n_398)
    | ((csa_tree_add_106_2_groupi_n_398 & csa_tree_add_106_2_groupi_n_705) | (csa_tree_add_106_2_groupi_n_705
    & csa_tree_add_106_2_groupi_n_788)));
 assign csa_tree_add_106_2_groupi_n_823 = (csa_tree_add_106_2_groupi_n_398 ^ (csa_tree_add_106_2_groupi_n_705
    ^ csa_tree_add_106_2_groupi_n_788));
 assign csa_tree_add_106_2_groupi_n_819 = ((csa_tree_add_106_2_groupi_n_782 & csa_tree_add_106_2_groupi_n_399)
    | ((csa_tree_add_106_2_groupi_n_399 & csa_tree_add_106_2_groupi_n_732) | (csa_tree_add_106_2_groupi_n_732
    & csa_tree_add_106_2_groupi_n_782)));
 assign csa_tree_add_106_2_groupi_n_820 = (csa_tree_add_106_2_groupi_n_399 ^ (csa_tree_add_106_2_groupi_n_732
    ^ csa_tree_add_106_2_groupi_n_782));
 assign csa_tree_add_106_2_groupi_n_817 = ((csa_tree_add_106_2_groupi_n_749 & csa_tree_add_106_2_groupi_n_748)
    | ((csa_tree_add_106_2_groupi_n_748 & csa_tree_add_106_2_groupi_n_699) | (csa_tree_add_106_2_groupi_n_699
    & csa_tree_add_106_2_groupi_n_749)));
 assign csa_tree_add_106_2_groupi_n_818 = (csa_tree_add_106_2_groupi_n_748 ^ (csa_tree_add_106_2_groupi_n_699
    ^ csa_tree_add_106_2_groupi_n_749));
 assign csa_tree_add_106_2_groupi_n_815 = ((csa_tree_add_106_2_groupi_n_752 & csa_tree_add_106_2_groupi_n_684)
    | ((csa_tree_add_106_2_groupi_n_684 & csa_tree_add_106_2_groupi_n_353) | (csa_tree_add_106_2_groupi_n_353
    & csa_tree_add_106_2_groupi_n_752)));
 assign csa_tree_add_106_2_groupi_n_816 = (csa_tree_add_106_2_groupi_n_684 ^ (csa_tree_add_106_2_groupi_n_353
    ^ csa_tree_add_106_2_groupi_n_752));
 assign csa_tree_add_106_2_groupi_n_813 = ((csa_tree_add_106_2_groupi_n_772 & csa_tree_add_106_2_groupi_n_397)
    | ((csa_tree_add_106_2_groupi_n_397 & csa_tree_add_106_2_groupi_n_730) | (csa_tree_add_106_2_groupi_n_730
    & csa_tree_add_106_2_groupi_n_772)));
 assign csa_tree_add_106_2_groupi_n_814 = (csa_tree_add_106_2_groupi_n_397 ^ (csa_tree_add_106_2_groupi_n_730
    ^ csa_tree_add_106_2_groupi_n_772));
 assign csa_tree_add_106_2_groupi_n_811 = ((csa_tree_add_106_2_groupi_n_774 & csa_tree_add_106_2_groupi_n_721)
    | ((csa_tree_add_106_2_groupi_n_721 & csa_tree_add_106_2_groupi_n_728) | (csa_tree_add_106_2_groupi_n_728
    & csa_tree_add_106_2_groupi_n_774)));
 assign csa_tree_add_106_2_groupi_n_812 = (csa_tree_add_106_2_groupi_n_721 ^ (csa_tree_add_106_2_groupi_n_728
    ^ csa_tree_add_106_2_groupi_n_774));
 assign csa_tree_add_106_2_groupi_n_809 = ((csa_tree_add_106_2_groupi_n_743 & csa_tree_add_106_2_groupi_n_386)
    | ((csa_tree_add_106_2_groupi_n_386 & csa_tree_add_106_2_groupi_n_711) | (csa_tree_add_106_2_groupi_n_711
    & csa_tree_add_106_2_groupi_n_743)));
 assign csa_tree_add_106_2_groupi_n_810 = (csa_tree_add_106_2_groupi_n_386 ^ (csa_tree_add_106_2_groupi_n_711
    ^ csa_tree_add_106_2_groupi_n_743));
 assign csa_tree_add_106_2_groupi_n_807 = ((csa_tree_add_106_2_groupi_n_780 & csa_tree_add_106_2_groupi_n_403)
    | ((csa_tree_add_106_2_groupi_n_403 & csa_tree_add_106_2_groupi_n_713) | (csa_tree_add_106_2_groupi_n_713
    & csa_tree_add_106_2_groupi_n_780)));
 assign csa_tree_add_106_2_groupi_n_808 = (csa_tree_add_106_2_groupi_n_403 ^ (csa_tree_add_106_2_groupi_n_713
    ^ csa_tree_add_106_2_groupi_n_780));
 assign csa_tree_add_106_2_groupi_n_805 = ((csa_tree_add_106_2_groupi_n_741 & csa_tree_add_106_2_groupi_n_411)
    | ((csa_tree_add_106_2_groupi_n_411 & csa_tree_add_106_2_groupi_n_720) | (csa_tree_add_106_2_groupi_n_720
    & csa_tree_add_106_2_groupi_n_741)));
 assign csa_tree_add_106_2_groupi_n_806 = (csa_tree_add_106_2_groupi_n_411 ^ (csa_tree_add_106_2_groupi_n_720
    ^ csa_tree_add_106_2_groupi_n_741));
 assign csa_tree_add_106_2_groupi_n_801 = ((csa_tree_add_106_2_groupi_n_768 & csa_tree_add_106_2_groupi_n_540)
    | ((csa_tree_add_106_2_groupi_n_540 & csa_tree_add_106_2_groupi_n_715) | (csa_tree_add_106_2_groupi_n_715
    & csa_tree_add_106_2_groupi_n_768)));
 assign csa_tree_add_106_2_groupi_n_802 = (csa_tree_add_106_2_groupi_n_540 ^ (csa_tree_add_106_2_groupi_n_715
    ^ csa_tree_add_106_2_groupi_n_768));
 assign csa_tree_add_106_2_groupi_n_795 = ((csa_tree_add_106_2_groupi_n_722 & csa_tree_add_106_2_groupi_n_387)
    | ((csa_tree_add_106_2_groupi_n_387 & csa_tree_add_106_2_groupi_n_723) | (csa_tree_add_106_2_groupi_n_723
    & csa_tree_add_106_2_groupi_n_722)));
 assign csa_tree_add_106_2_groupi_n_796 = (csa_tree_add_106_2_groupi_n_387 ^ (csa_tree_add_106_2_groupi_n_723
    ^ csa_tree_add_106_2_groupi_n_722));
 assign csa_tree_add_106_2_groupi_n_791 = ((csa_tree_add_106_2_groupi_n_757 & csa_tree_add_106_2_groupi_n_544)
    | ((csa_tree_add_106_2_groupi_n_544 & csa_tree_add_106_2_groupi_n_691) | (csa_tree_add_106_2_groupi_n_691
    & csa_tree_add_106_2_groupi_n_757)));
 assign csa_tree_add_106_2_groupi_n_792 = (csa_tree_add_106_2_groupi_n_544 ^ (csa_tree_add_106_2_groupi_n_691
    ^ csa_tree_add_106_2_groupi_n_757));
 assign csa_tree_add_106_2_groupi_n_788 = ((csa_tree_add_106_2_groupi_n_753 & csa_tree_add_106_2_groupi_n_600)
    | ((csa_tree_add_106_2_groupi_n_600 & csa_tree_add_106_2_groupi_n_657) | (csa_tree_add_106_2_groupi_n_657
    & csa_tree_add_106_2_groupi_n_753)));
 assign csa_tree_add_106_2_groupi_n_789 = (csa_tree_add_106_2_groupi_n_600 ^ (csa_tree_add_106_2_groupi_n_657
    ^ csa_tree_add_106_2_groupi_n_753));
 assign csa_tree_add_106_2_groupi_n_786 = ((csa_tree_add_106_2_groupi_n_751 & csa_tree_add_106_2_groupi_n_589)
    | ((csa_tree_add_106_2_groupi_n_589 & csa_tree_add_106_2_groupi_n_472) | (csa_tree_add_106_2_groupi_n_472
    & csa_tree_add_106_2_groupi_n_751)));
 assign csa_tree_add_106_2_groupi_n_787 = (csa_tree_add_106_2_groupi_n_589 ^ (csa_tree_add_106_2_groupi_n_472
    ^ csa_tree_add_106_2_groupi_n_751));
 assign csa_tree_add_106_2_groupi_n_784 = ((csa_tree_add_106_2_groupi_n_733 & csa_tree_add_106_2_groupi_n_542)
    | ((csa_tree_add_106_2_groupi_n_542 & csa_tree_add_106_2_groupi_n_709) | (csa_tree_add_106_2_groupi_n_709
    & csa_tree_add_106_2_groupi_n_733)));
 assign csa_tree_add_106_2_groupi_n_785 = (csa_tree_add_106_2_groupi_n_542 ^ (csa_tree_add_106_2_groupi_n_709
    ^ csa_tree_add_106_2_groupi_n_733));
 assign csa_tree_add_106_2_groupi_n_782 = ((csa_tree_add_106_2_groupi_n_729 & csa_tree_add_106_2_groupi_n_571)
    | ((csa_tree_add_106_2_groupi_n_571 & csa_tree_add_106_2_groupi_n_479) | (csa_tree_add_106_2_groupi_n_479
    & csa_tree_add_106_2_groupi_n_729)));
 assign csa_tree_add_106_2_groupi_n_783 = (csa_tree_add_106_2_groupi_n_571 ^ (csa_tree_add_106_2_groupi_n_479
    ^ csa_tree_add_106_2_groupi_n_729));
 assign csa_tree_add_106_2_groupi_n_780 = ((csa_tree_add_106_2_groupi_n_731 & csa_tree_add_106_2_groupi_n_547)
    | ((csa_tree_add_106_2_groupi_n_547 & csa_tree_add_106_2_groupi_n_671) | (csa_tree_add_106_2_groupi_n_671
    & csa_tree_add_106_2_groupi_n_731)));
 assign csa_tree_add_106_2_groupi_n_781 = (csa_tree_add_106_2_groupi_n_547 ^ (csa_tree_add_106_2_groupi_n_671
    ^ csa_tree_add_106_2_groupi_n_731));
 assign csa_tree_add_106_2_groupi_n_778 = ((csa_tree_add_106_2_groupi_n_707 & csa_tree_add_106_2_groupi_n_496)
    | ((csa_tree_add_106_2_groupi_n_496 & csa_tree_add_106_2_groupi_n_491) | (csa_tree_add_106_2_groupi_n_491
    & csa_tree_add_106_2_groupi_n_707)));
 assign csa_tree_add_106_2_groupi_n_779 = (csa_tree_add_106_2_groupi_n_496 ^ (csa_tree_add_106_2_groupi_n_491
    ^ csa_tree_add_106_2_groupi_n_707));
 assign csa_tree_add_106_2_groupi_n_776 = ((csa_tree_add_106_2_groupi_n_719 & csa_tree_add_106_2_groupi_n_652)
    | ((csa_tree_add_106_2_groupi_n_652 & csa_tree_add_106_2_groupi_n_673) | (csa_tree_add_106_2_groupi_n_673
    & csa_tree_add_106_2_groupi_n_719)));
 assign csa_tree_add_106_2_groupi_n_777 = (csa_tree_add_106_2_groupi_n_652 ^ (csa_tree_add_106_2_groupi_n_673
    ^ csa_tree_add_106_2_groupi_n_719));
 assign csa_tree_add_106_2_groupi_n_774 = ((csa_tree_add_106_2_groupi_n_708 & csa_tree_add_106_2_groupi_n_601)
    | ((csa_tree_add_106_2_groupi_n_601 & csa_tree_add_106_2_groupi_n_475) | (csa_tree_add_106_2_groupi_n_475
    & csa_tree_add_106_2_groupi_n_708)));
 assign csa_tree_add_106_2_groupi_n_775 = (csa_tree_add_106_2_groupi_n_601 ^ (csa_tree_add_106_2_groupi_n_475
    ^ csa_tree_add_106_2_groupi_n_708));
 assign csa_tree_add_106_2_groupi_n_772 = ((csa_tree_add_106_2_groupi_n_727 & csa_tree_add_106_2_groupi_n_564)
    | ((csa_tree_add_106_2_groupi_n_564 & csa_tree_add_106_2_groupi_n_468) | (csa_tree_add_106_2_groupi_n_468
    & csa_tree_add_106_2_groupi_n_727)));
 assign csa_tree_add_106_2_groupi_n_773 = (csa_tree_add_106_2_groupi_n_564 ^ (csa_tree_add_106_2_groupi_n_468
    ^ csa_tree_add_106_2_groupi_n_727));
 assign csa_tree_add_106_2_groupi_n_770 = ((csa_tree_add_106_2_groupi_n_706 & csa_tree_add_106_2_groupi_n_503)
    | ((csa_tree_add_106_2_groupi_n_503 & csa_tree_add_106_2_groupi_n_639) | (csa_tree_add_106_2_groupi_n_639
    & csa_tree_add_106_2_groupi_n_706)));
 assign csa_tree_add_106_2_groupi_n_771 = (csa_tree_add_106_2_groupi_n_503 ^ (csa_tree_add_106_2_groupi_n_639
    ^ csa_tree_add_106_2_groupi_n_706));
 assign csa_tree_add_106_2_groupi_n_768 = ((csa_tree_add_106_2_groupi_n_702 & csa_tree_add_106_2_groupi_n_478)
    | ((csa_tree_add_106_2_groupi_n_478 & csa_tree_add_106_2_groupi_n_523) | (csa_tree_add_106_2_groupi_n_523
    & csa_tree_add_106_2_groupi_n_702)));
 assign csa_tree_add_106_2_groupi_n_769 = (csa_tree_add_106_2_groupi_n_478 ^ (csa_tree_add_106_2_groupi_n_523
    ^ csa_tree_add_106_2_groupi_n_702));
 assign csa_tree_add_106_2_groupi_n_767 = ~(csa_tree_add_106_2_groupi_n_739 ^ csa_tree_add_106_2_groupi_n_674);
 assign csa_tree_add_106_2_groupi_n_763 = ((csa_tree_add_106_2_groupi_n_703 & csa_tree_add_106_2_groupi_n_514)
    | ((csa_tree_add_106_2_groupi_n_514 & csa_tree_add_106_2_groupi_n_675) | (csa_tree_add_106_2_groupi_n_675
    & csa_tree_add_106_2_groupi_n_703)));
 assign csa_tree_add_106_2_groupi_n_764 = (csa_tree_add_106_2_groupi_n_514 ^ (csa_tree_add_106_2_groupi_n_675
    ^ csa_tree_add_106_2_groupi_n_703));
 assign csa_tree_add_106_2_groupi_n_761 = ((csa_tree_add_106_2_groupi_n_697 & csa_tree_add_106_2_groupi_n_455)
    | ((csa_tree_add_106_2_groupi_n_455 & csa_tree_add_106_2_groupi_n_463) | (csa_tree_add_106_2_groupi_n_463
    & csa_tree_add_106_2_groupi_n_697)));
 assign csa_tree_add_106_2_groupi_n_762 = (csa_tree_add_106_2_groupi_n_455 ^ (csa_tree_add_106_2_groupi_n_463
    ^ csa_tree_add_106_2_groupi_n_697));
 assign csa_tree_add_106_2_groupi_n_757 = ((csa_tree_add_106_2_groupi_n_678 & csa_tree_add_106_2_groupi_n_481)
    | ((csa_tree_add_106_2_groupi_n_481 & csa_tree_add_106_2_groupi_n_402) | (csa_tree_add_106_2_groupi_n_402
    & csa_tree_add_106_2_groupi_n_678)));
 assign csa_tree_add_106_2_groupi_n_758 = (csa_tree_add_106_2_groupi_n_481 ^ (csa_tree_add_106_2_groupi_n_402
    ^ csa_tree_add_106_2_groupi_n_678));
 assign csa_tree_add_106_2_groupi_n_753 = ((csa_tree_add_106_2_groupi_n_659 & csa_tree_add_106_2_groupi_n_520)
    | ((csa_tree_add_106_2_groupi_n_520 & csa_tree_add_106_2_groupi_n_666) | (csa_tree_add_106_2_groupi_n_666
    & csa_tree_add_106_2_groupi_n_659)));
 assign csa_tree_add_106_2_groupi_n_754 = (csa_tree_add_106_2_groupi_n_520 ^ (csa_tree_add_106_2_groupi_n_666
    ^ csa_tree_add_106_2_groupi_n_659));
 assign csa_tree_add_106_2_groupi_n_751 = ((csa_tree_add_106_2_groupi_n_663 & csa_tree_add_106_2_groupi_n_516)
    | ((csa_tree_add_106_2_groupi_n_516 & csa_tree_add_106_2_groupi_n_654) | (csa_tree_add_106_2_groupi_n_654
    & csa_tree_add_106_2_groupi_n_663)));
 assign csa_tree_add_106_2_groupi_n_752 = (csa_tree_add_106_2_groupi_n_516 ^ (csa_tree_add_106_2_groupi_n_654
    ^ csa_tree_add_106_2_groupi_n_663));
 assign csa_tree_add_106_2_groupi_n_749 = ((csa_tree_add_106_2_groupi_n_700 & csa_tree_add_106_2_groupi_n_672)
    | ((csa_tree_add_106_2_groupi_n_672 & csa_tree_add_106_2_groupi_n_643) | (csa_tree_add_106_2_groupi_n_643
    & csa_tree_add_106_2_groupi_n_700)));
 assign csa_tree_add_106_2_groupi_n_750 = (csa_tree_add_106_2_groupi_n_672 ^ (csa_tree_add_106_2_groupi_n_643
    ^ csa_tree_add_106_2_groupi_n_700));
 assign csa_tree_add_106_2_groupi_n_747 = ((csa_tree_add_106_2_groupi_n_688 & csa_tree_add_106_2_groupi_n_642)
    | ((csa_tree_add_106_2_groupi_n_642 & csa_tree_add_106_2_groupi_n_669) | (csa_tree_add_106_2_groupi_n_669
    & csa_tree_add_106_2_groupi_n_688)));
 assign csa_tree_add_106_2_groupi_n_748 = (csa_tree_add_106_2_groupi_n_642 ^ (csa_tree_add_106_2_groupi_n_669
    ^ csa_tree_add_106_2_groupi_n_688));
 assign csa_tree_add_106_2_groupi_n_745 = ((csa_tree_add_106_2_groupi_n_676 & csa_tree_add_106_2_groupi_n_476)
    | ((csa_tree_add_106_2_groupi_n_476 & csa_tree_add_106_2_groupi_n_551) | (csa_tree_add_106_2_groupi_n_551
    & csa_tree_add_106_2_groupi_n_676)));
 assign csa_tree_add_106_2_groupi_n_746 = (csa_tree_add_106_2_groupi_n_476 ^ (csa_tree_add_106_2_groupi_n_551
    ^ csa_tree_add_106_2_groupi_n_676));
 assign csa_tree_add_106_2_groupi_n_743 = ((csa_tree_add_106_2_groupi_n_704 & csa_tree_add_106_2_groupi_n_670)
    | ((csa_tree_add_106_2_groupi_n_670 & csa_tree_add_106_2_groupi_n_485) | (csa_tree_add_106_2_groupi_n_485
    & csa_tree_add_106_2_groupi_n_704)));
 assign csa_tree_add_106_2_groupi_n_744 = (csa_tree_add_106_2_groupi_n_670 ^ (csa_tree_add_106_2_groupi_n_485
    ^ csa_tree_add_106_2_groupi_n_704));
 assign csa_tree_add_106_2_groupi_n_741 = ((csa_tree_add_106_2_groupi_n_712 & csa_tree_add_106_2_groupi_n_471)
    | ((csa_tree_add_106_2_groupi_n_471 & csa_tree_add_106_2_groupi_n_650) | (csa_tree_add_106_2_groupi_n_650
    & csa_tree_add_106_2_groupi_n_712)));
 assign csa_tree_add_106_2_groupi_n_742 = (csa_tree_add_106_2_groupi_n_471 ^ (csa_tree_add_106_2_groupi_n_650
    ^ csa_tree_add_106_2_groupi_n_712));
 assign csa_tree_add_106_2_groupi_n_739 = ((csa_tree_add_106_2_groupi_n_682 & csa_tree_add_106_2_groupi_n_644)
    | ((csa_tree_add_106_2_groupi_n_644 & csa_tree_add_106_2_groupi_n_641) | (csa_tree_add_106_2_groupi_n_641
    & csa_tree_add_106_2_groupi_n_682)));
 assign csa_tree_add_106_2_groupi_n_740 = (csa_tree_add_106_2_groupi_n_644 ^ (csa_tree_add_106_2_groupi_n_641
    ^ csa_tree_add_106_2_groupi_n_682));
 assign csa_tree_add_106_2_groupi_n_737 = ((csa_tree_add_106_2_groupi_n_710 & csa_tree_add_106_2_groupi_n_582)
    | ((csa_tree_add_106_2_groupi_n_582 & csa_tree_add_106_2_groupi_n_653) | (csa_tree_add_106_2_groupi_n_653
    & csa_tree_add_106_2_groupi_n_710)));
 assign csa_tree_add_106_2_groupi_n_738 = (csa_tree_add_106_2_groupi_n_582 ^ (csa_tree_add_106_2_groupi_n_653
    ^ csa_tree_add_106_2_groupi_n_710));
 assign csa_tree_add_106_2_groupi_n_735 = ((csa_tree_add_106_2_groupi_n_698 & csa_tree_add_106_2_groupi_n_668)
    | ((csa_tree_add_106_2_groupi_n_668 & csa_tree_add_106_2_groupi_n_645) | (csa_tree_add_106_2_groupi_n_645
    & csa_tree_add_106_2_groupi_n_698)));
 assign csa_tree_add_106_2_groupi_n_736 = (csa_tree_add_106_2_groupi_n_668 ^ (csa_tree_add_106_2_groupi_n_645
    ^ csa_tree_add_106_2_groupi_n_698));
 assign csa_tree_add_106_2_groupi_n_733 = ((csa_tree_add_106_2_groupi_n_714 & csa_tree_add_106_2_groupi_n_482)
    | ((csa_tree_add_106_2_groupi_n_482 & csa_tree_add_106_2_groupi_n_409) | (csa_tree_add_106_2_groupi_n_409
    & csa_tree_add_106_2_groupi_n_714)));
 assign csa_tree_add_106_2_groupi_n_734 = (csa_tree_add_106_2_groupi_n_482 ^ (csa_tree_add_106_2_groupi_n_409
    ^ csa_tree_add_106_2_groupi_n_714));
 assign csa_tree_add_106_2_groupi_n_731 = ((csa_tree_add_106_2_groupi_n_658 & csa_tree_add_106_2_groupi_n_480)
    | ((csa_tree_add_106_2_groupi_n_480 & csa_tree_add_106_2_groupi_n_526) | (csa_tree_add_106_2_groupi_n_526
    & csa_tree_add_106_2_groupi_n_658)));
 assign csa_tree_add_106_2_groupi_n_732 = (csa_tree_add_106_2_groupi_n_480 ^ (csa_tree_add_106_2_groupi_n_526
    ^ csa_tree_add_106_2_groupi_n_658));
 assign csa_tree_add_106_2_groupi_n_729 = ((csa_tree_add_106_2_groupi_n_667 & csa_tree_add_106_2_groupi_n_511)
    | ((csa_tree_add_106_2_groupi_n_511 & csa_tree_add_106_2_groupi_n_662) | (csa_tree_add_106_2_groupi_n_662
    & csa_tree_add_106_2_groupi_n_667)));
 assign csa_tree_add_106_2_groupi_n_730 = (csa_tree_add_106_2_groupi_n_511 ^ (csa_tree_add_106_2_groupi_n_662
    ^ csa_tree_add_106_2_groupi_n_667));
 assign csa_tree_add_106_2_groupi_n_727 = ((csa_tree_add_106_2_groupi_n_648 & csa_tree_add_106_2_groupi_n_494)
    | ((csa_tree_add_106_2_groupi_n_494 & csa_tree_add_106_2_groupi_n_655) | (csa_tree_add_106_2_groupi_n_655
    & csa_tree_add_106_2_groupi_n_648)));
 assign csa_tree_add_106_2_groupi_n_728 = (csa_tree_add_106_2_groupi_n_494 ^ (csa_tree_add_106_2_groupi_n_655
    ^ csa_tree_add_106_2_groupi_n_648));
 assign csa_tree_add_106_2_groupi_n_723 = ((csa_tree_add_106_2_groupi_n_690 & csa_tree_add_106_2_groupi_n_389)
    | ((csa_tree_add_106_2_groupi_n_389 & csa_tree_add_106_2_groupi_n_461) | (csa_tree_add_106_2_groupi_n_461
    & csa_tree_add_106_2_groupi_n_690)));
 assign csa_tree_add_106_2_groupi_n_724 = (csa_tree_add_106_2_groupi_n_389 ^ (csa_tree_add_106_2_groupi_n_461
    ^ csa_tree_add_106_2_groupi_n_690));
 assign csa_tree_add_106_2_groupi_n_721 = ((csa_tree_add_106_2_groupi_n_649 & csa_tree_add_106_2_groupi_n_486)
    | ((csa_tree_add_106_2_groupi_n_486 & csa_tree_add_106_2_groupi_n_646) | (csa_tree_add_106_2_groupi_n_646
    & csa_tree_add_106_2_groupi_n_649)));
 assign csa_tree_add_106_2_groupi_n_722 = (csa_tree_add_106_2_groupi_n_486 ^ (csa_tree_add_106_2_groupi_n_646
    ^ csa_tree_add_106_2_groupi_n_649));
 assign csa_tree_add_106_2_groupi_n_719 = ((csa_tree_add_106_2_groupi_n_664 & csa_tree_add_106_2_groupi_n_467)
    | ((csa_tree_add_106_2_groupi_n_467 & csa_tree_add_106_2_groupi_n_495) | (csa_tree_add_106_2_groupi_n_495
    & csa_tree_add_106_2_groupi_n_664)));
 assign csa_tree_add_106_2_groupi_n_720 = (csa_tree_add_106_2_groupi_n_467 ^ (csa_tree_add_106_2_groupi_n_495
    ^ csa_tree_add_106_2_groupi_n_664));
 assign csa_tree_add_106_2_groupi_n_717 = ((csa_tree_add_106_2_groupi_n_660 & csa_tree_add_106_2_groupi_n_592)
    | ((csa_tree_add_106_2_groupi_n_592 & csa_tree_add_106_2_groupi_n_635) | (csa_tree_add_106_2_groupi_n_635
    & csa_tree_add_106_2_groupi_n_660)));
 assign csa_tree_add_106_2_groupi_n_718 = (csa_tree_add_106_2_groupi_n_592 ^ (csa_tree_add_106_2_groupi_n_635
    ^ csa_tree_add_106_2_groupi_n_660));
 assign csa_tree_add_106_2_groupi_n_716 = ~(csa_tree_add_106_2_groupi_n_680 ^ csa_tree_add_106_2_groupi_n_677);
 assign csa_tree_add_106_2_groupi_n_714 = ((csa_tree_add_106_2_groupi_n_532 & csa_tree_add_106_2_groupi_n_581)
    | ((csa_tree_add_106_2_groupi_n_581 & csa_tree_add_106_2_groupi_n_408) | (csa_tree_add_106_2_groupi_n_408
    & csa_tree_add_106_2_groupi_n_532)));
 assign csa_tree_add_106_2_groupi_n_715 = (csa_tree_add_106_2_groupi_n_581 ^ (csa_tree_add_106_2_groupi_n_408
    ^ csa_tree_add_106_2_groupi_n_532));
 assign csa_tree_add_106_2_groupi_n_712 = ((csa_tree_add_106_2_groupi_n_651 & csa_tree_add_106_2_groupi_n_596)
    | ((csa_tree_add_106_2_groupi_n_596 & csa_tree_add_106_2_groupi_n_501) | (csa_tree_add_106_2_groupi_n_501
    & csa_tree_add_106_2_groupi_n_651)));
 assign csa_tree_add_106_2_groupi_n_713 = (csa_tree_add_106_2_groupi_n_596 ^ (csa_tree_add_106_2_groupi_n_501
    ^ csa_tree_add_106_2_groupi_n_651));
 assign csa_tree_add_106_2_groupi_n_710 = ((csa_tree_add_106_2_groupi_n_665 & csa_tree_add_106_2_groupi_n_585)
    | ((csa_tree_add_106_2_groupi_n_585 & csa_tree_add_106_2_groupi_n_508) | (csa_tree_add_106_2_groupi_n_508
    & csa_tree_add_106_2_groupi_n_665)));
 assign csa_tree_add_106_2_groupi_n_711 = (csa_tree_add_106_2_groupi_n_585 ^ (csa_tree_add_106_2_groupi_n_508
    ^ csa_tree_add_106_2_groupi_n_665));
 assign csa_tree_add_106_2_groupi_n_708 = (csa_tree_add_106_2_groupi_n_647 & csa_tree_add_106_2_groupi_n_529);
 assign csa_tree_add_106_2_groupi_n_709 = (csa_tree_add_106_2_groupi_n_647 ^ csa_tree_add_106_2_groupi_n_529);
 assign csa_tree_add_106_2_groupi_n_706 = ((csa_tree_add_106_2_groupi_n_636 & csa_tree_add_106_2_groupi_n_536)
    | ((csa_tree_add_106_2_groupi_n_536 & csa_tree_add_106_2_groupi_n_534) | (csa_tree_add_106_2_groupi_n_534
    & csa_tree_add_106_2_groupi_n_636)));
 assign csa_tree_add_106_2_groupi_n_707 = (csa_tree_add_106_2_groupi_n_536 ^ (csa_tree_add_106_2_groupi_n_534
    ^ csa_tree_add_106_2_groupi_n_636));
 assign csa_tree_add_106_2_groupi_n_704 = ((csa_tree_add_106_2_groupi_n_656 & csa_tree_add_106_2_groupi_n_460)
    | ((csa_tree_add_106_2_groupi_n_460 & csa_tree_add_106_2_groupi_n_579) | (csa_tree_add_106_2_groupi_n_579
    & csa_tree_add_106_2_groupi_n_656)));
 assign csa_tree_add_106_2_groupi_n_705 = (csa_tree_add_106_2_groupi_n_460 ^ (csa_tree_add_106_2_groupi_n_579
    ^ csa_tree_add_106_2_groupi_n_656));
 assign csa_tree_add_106_2_groupi_n_702 = ((csa_tree_add_106_2_groupi_n_422 & csa_tree_add_106_2_groupi_n_570)
    | ((csa_tree_add_106_2_groupi_n_570 & csa_tree_add_106_2_groupi_n_404) | (csa_tree_add_106_2_groupi_n_404
    & csa_tree_add_106_2_groupi_n_422)));
 assign csa_tree_add_106_2_groupi_n_703 = (csa_tree_add_106_2_groupi_n_570 ^ (csa_tree_add_106_2_groupi_n_404
    ^ csa_tree_add_106_2_groupi_n_422));
 assign csa_tree_add_106_2_groupi_n_700 = ((csa_tree_add_106_2_groupi_n_608 & csa_tree_add_106_2_groupi_n_528)
    | ((csa_tree_add_106_2_groupi_n_528 & csa_tree_add_106_2_groupi_n_483) | (csa_tree_add_106_2_groupi_n_483
    & csa_tree_add_106_2_groupi_n_608)));
 assign csa_tree_add_106_2_groupi_n_701 = (csa_tree_add_106_2_groupi_n_528 ^ (csa_tree_add_106_2_groupi_n_483
    ^ csa_tree_add_106_2_groupi_n_608));
 assign csa_tree_add_106_2_groupi_n_698 = ((csa_tree_add_106_2_groupi_n_610 & csa_tree_add_106_2_groupi_n_586)
    | ((csa_tree_add_106_2_groupi_n_586 & csa_tree_add_106_2_groupi_n_572) | (csa_tree_add_106_2_groupi_n_572
    & csa_tree_add_106_2_groupi_n_610)));
 assign csa_tree_add_106_2_groupi_n_699 = (csa_tree_add_106_2_groupi_n_586 ^ (csa_tree_add_106_2_groupi_n_572
    ^ csa_tree_add_106_2_groupi_n_610));
 assign csa_tree_add_106_2_groupi_n_696 = ((csa_tree_add_106_2_groupi_n_605 & csa_tree_add_106_2_groupi_n_538)
    | ((csa_tree_add_106_2_groupi_n_538 & csa_tree_add_106_2_groupi_n_634) | (csa_tree_add_106_2_groupi_n_634
    & csa_tree_add_106_2_groupi_n_605)));
 assign csa_tree_add_106_2_groupi_n_697 = (csa_tree_add_106_2_groupi_n_538 ^ (csa_tree_add_106_2_groupi_n_634
    ^ csa_tree_add_106_2_groupi_n_605));
 assign csa_tree_add_106_2_groupi_n_690 = ((csa_tree_add_106_2_groupi_n_615 & csa_tree_add_106_2_groupi_n_535)
    | ((csa_tree_add_106_2_groupi_n_535 & csa_tree_add_106_2_groupi_n_401) | (csa_tree_add_106_2_groupi_n_401
    & csa_tree_add_106_2_groupi_n_615)));
 assign csa_tree_add_106_2_groupi_n_691 = (csa_tree_add_106_2_groupi_n_535 ^ (csa_tree_add_106_2_groupi_n_401
    ^ csa_tree_add_106_2_groupi_n_615));
 assign csa_tree_add_106_2_groupi_n_688 = ((csa_tree_add_106_2_groupi_n_625 & csa_tree_add_106_2_groupi_n_587)
    | ((csa_tree_add_106_2_groupi_n_587 & csa_tree_add_106_2_groupi_n_470) | (csa_tree_add_106_2_groupi_n_470
    & csa_tree_add_106_2_groupi_n_625)));
 assign csa_tree_add_106_2_groupi_n_689 = (csa_tree_add_106_2_groupi_n_587 ^ (csa_tree_add_106_2_groupi_n_470
    ^ csa_tree_add_106_2_groupi_n_625));
 assign csa_tree_add_106_2_groupi_n_686 = ((csa_tree_add_106_2_groupi_n_617 & csa_tree_add_106_2_groupi_n_638)
    | ((csa_tree_add_106_2_groupi_n_638 & csa_tree_add_106_2_groupi_n_584) | (csa_tree_add_106_2_groupi_n_584
    & csa_tree_add_106_2_groupi_n_617)));
 assign csa_tree_add_106_2_groupi_n_687 = (csa_tree_add_106_2_groupi_n_638 ^ (csa_tree_add_106_2_groupi_n_584
    ^ csa_tree_add_106_2_groupi_n_617));
 assign csa_tree_add_106_2_groupi_n_684 = ((csa_tree_add_106_2_groupi_n_612 & csa_tree_add_106_2_groupi_n_395)
    | ((csa_tree_add_106_2_groupi_n_395 & csa_tree_add_106_2_groupi_n_464) | (csa_tree_add_106_2_groupi_n_464
    & csa_tree_add_106_2_groupi_n_612)));
 assign csa_tree_add_106_2_groupi_n_685 = (csa_tree_add_106_2_groupi_n_395 ^ (csa_tree_add_106_2_groupi_n_464
    ^ csa_tree_add_106_2_groupi_n_612));
 assign csa_tree_add_106_2_groupi_n_682 = ((csa_tree_add_106_2_groupi_n_606 & csa_tree_add_106_2_groupi_n_539)
    | ((csa_tree_add_106_2_groupi_n_539 & csa_tree_add_106_2_groupi_n_513) | (csa_tree_add_106_2_groupi_n_513
    & csa_tree_add_106_2_groupi_n_606)));
 assign csa_tree_add_106_2_groupi_n_683 = (csa_tree_add_106_2_groupi_n_539 ^ (csa_tree_add_106_2_groupi_n_513
    ^ csa_tree_add_106_2_groupi_n_606));
 assign csa_tree_add_106_2_groupi_n_680 = ((csa_tree_add_106_2_groupi_n_609 & csa_tree_add_106_2_groupi_n_598)
    | ((csa_tree_add_106_2_groupi_n_598 & csa_tree_add_106_2_groupi_n_575) | (csa_tree_add_106_2_groupi_n_575
    & csa_tree_add_106_2_groupi_n_609)));
 assign csa_tree_add_106_2_groupi_n_681 = (csa_tree_add_106_2_groupi_n_598 ^ (csa_tree_add_106_2_groupi_n_575
    ^ csa_tree_add_106_2_groupi_n_609));
 assign csa_tree_add_106_2_groupi_n_678 = ((csa_tree_add_106_2_groupi_n_417 & csa_tree_add_106_2_groupi_n_577)
    | ((csa_tree_add_106_2_groupi_n_577 & csa_tree_add_106_2_groupi_n_405) | (csa_tree_add_106_2_groupi_n_405
    & csa_tree_add_106_2_groupi_n_417)));
 assign csa_tree_add_106_2_groupi_n_679 = (csa_tree_add_106_2_groupi_n_577 ^ (csa_tree_add_106_2_groupi_n_405
    ^ csa_tree_add_106_2_groupi_n_417));
 assign csa_tree_add_106_2_groupi_n_677 = ~(csa_tree_add_106_2_groupi_n_633 ^ csa_tree_add_106_2_groupi_n_426);
 assign csa_tree_add_106_2_groupi_n_674 = ~(csa_tree_add_106_2_groupi_n_640 ^ csa_tree_add_106_2_groupi_n_626);
 assign csa_tree_add_106_2_groupi_n_672 = (csa_tree_add_106_2_groupi_n_623 & csa_tree_add_106_2_groupi_n_413);
 assign csa_tree_add_106_2_groupi_n_673 = (csa_tree_add_106_2_groupi_n_623 ^ csa_tree_add_106_2_groupi_n_413);
 assign csa_tree_add_106_2_groupi_n_670 = (csa_tree_add_106_2_groupi_n_530 & csa_tree_add_106_2_groupi_n_416);
 assign csa_tree_add_106_2_groupi_n_671 = (csa_tree_add_106_2_groupi_n_530 ^ csa_tree_add_106_2_groupi_n_416);
 assign csa_tree_add_106_2_groupi_n_668 = (csa_tree_add_106_2_groupi_n_531 & csa_tree_add_106_2_groupi_n_391);
 assign csa_tree_add_106_2_groupi_n_669 = (csa_tree_add_106_2_groupi_n_531 ^ csa_tree_add_106_2_groupi_n_391);
 assign csa_tree_add_106_2_groupi_n_666 = (csa_tree_add_106_2_groupi_n_619 & csa_tree_add_106_2_groupi_n_421);
 assign csa_tree_add_106_2_groupi_n_667 = (csa_tree_add_106_2_groupi_n_619 ^ csa_tree_add_106_2_groupi_n_421);
 assign csa_tree_add_106_2_groupi_n_664 = (csa_tree_add_106_2_groupi_n_607 & csa_tree_add_106_2_groupi_n_392);
 assign csa_tree_add_106_2_groupi_n_665 = (csa_tree_add_106_2_groupi_n_607 ^ csa_tree_add_106_2_groupi_n_392);
 assign csa_tree_add_106_2_groupi_n_662 = (csa_tree_add_106_2_groupi_n_620 & csa_tree_add_106_2_groupi_n_418);
 assign csa_tree_add_106_2_groupi_n_663 = (csa_tree_add_106_2_groupi_n_620 ^ csa_tree_add_106_2_groupi_n_418);
 assign csa_tree_add_106_2_groupi_n_660 = ((csa_tree_add_106_2_groupi_n_603 & csa_tree_add_106_2_groupi_n_207)
    | ((csa_tree_add_106_2_groupi_n_207 & csa_tree_add_106_2_groupi_n_208) | (csa_tree_add_106_2_groupi_n_208
    & csa_tree_add_106_2_groupi_n_603)));
 assign csa_tree_add_106_2_groupi_n_661 = (csa_tree_add_106_2_groupi_n_207 ^ (csa_tree_add_106_2_groupi_n_208
    ^ csa_tree_add_106_2_groupi_n_603));
 assign csa_tree_add_106_2_groupi_n_658 = (csa_tree_add_106_2_groupi_n_616 & csa_tree_add_106_2_groupi_n_412);
 assign csa_tree_add_106_2_groupi_n_659 = (csa_tree_add_106_2_groupi_n_616 ^ csa_tree_add_106_2_groupi_n_412);
 assign csa_tree_add_106_2_groupi_n_656 = (csa_tree_add_106_2_groupi_n_614 & csa_tree_add_106_2_groupi_n_414);
 assign csa_tree_add_106_2_groupi_n_657 = (csa_tree_add_106_2_groupi_n_614 ^ csa_tree_add_106_2_groupi_n_414);
 assign csa_tree_add_106_2_groupi_n_654 = (csa_tree_add_106_2_groupi_n_622 & csa_tree_add_106_2_groupi_n_424);
 assign csa_tree_add_106_2_groupi_n_655 = (csa_tree_add_106_2_groupi_n_622 ^ csa_tree_add_106_2_groupi_n_424);
 assign csa_tree_add_106_2_groupi_n_652 = (csa_tree_add_106_2_groupi_n_621 & csa_tree_add_106_2_groupi_n_415);
 assign csa_tree_add_106_2_groupi_n_653 = (csa_tree_add_106_2_groupi_n_621 ^ csa_tree_add_106_2_groupi_n_415);
 assign csa_tree_add_106_2_groupi_n_650 = (csa_tree_add_106_2_groupi_n_624 & csa_tree_add_106_2_groupi_n_390);
 assign csa_tree_add_106_2_groupi_n_651 = (csa_tree_add_106_2_groupi_n_624 ^ csa_tree_add_106_2_groupi_n_390);
 assign csa_tree_add_106_2_groupi_n_648 = (csa_tree_add_106_2_groupi_n_604 & csa_tree_add_106_2_groupi_n_425);
 assign csa_tree_add_106_2_groupi_n_649 = (csa_tree_add_106_2_groupi_n_604 ^ csa_tree_add_106_2_groupi_n_425);
 assign csa_tree_add_106_2_groupi_n_646 = (csa_tree_add_106_2_groupi_n_613 & csa_tree_add_106_2_groupi_n_393);
 assign csa_tree_add_106_2_groupi_n_647 = (csa_tree_add_106_2_groupi_n_613 ^ csa_tree_add_106_2_groupi_n_393);
 assign csa_tree_add_106_2_groupi_n_644 = (csa_tree_add_106_2_groupi_n_618 & csa_tree_add_106_2_groupi_n_423);
 assign csa_tree_add_106_2_groupi_n_645 = (csa_tree_add_106_2_groupi_n_618 ^ csa_tree_add_106_2_groupi_n_423);
 assign csa_tree_add_106_2_groupi_n_642 = (csa_tree_add_106_2_groupi_n_533 & csa_tree_add_106_2_groupi_n_420);
 assign csa_tree_add_106_2_groupi_n_643 = (csa_tree_add_106_2_groupi_n_533 ^ csa_tree_add_106_2_groupi_n_420);
 assign csa_tree_add_106_2_groupi_n_641 = ~(csa_tree_add_106_2_groupi_n_633 & (csa_tree_add_106_2_groupi_n_434
    | csa_tree_add_106_2_groupi_n_632));
 assign csa_tree_add_106_2_groupi_n_640 = ~(csa_tree_add_106_2_groupi_n_628 ^ csa_tree_add_106_2_groupi_n_5);
 assign csa_tree_add_106_2_groupi_n_638 = (csa_tree_add_106_2_groupi_n_349 & csa_tree_add_106_2_groupi_n_350);
 assign csa_tree_add_106_2_groupi_n_639 = (csa_tree_add_106_2_groupi_n_349 ^ csa_tree_add_106_2_groupi_n_350);
 assign csa_tree_add_106_2_groupi_n_636 = (csa_tree_add_106_2_groupi_n_347 & csa_tree_add_106_2_groupi_n_348);
 assign csa_tree_add_106_2_groupi_n_637 = (csa_tree_add_106_2_groupi_n_347 ^ csa_tree_add_106_2_groupi_n_348);
 assign csa_tree_add_106_2_groupi_n_634 = (csa_tree_add_106_2_groupi_n_346 & csa_tree_add_106_2_groupi_n_345);
 assign csa_tree_add_106_2_groupi_n_635 = (csa_tree_add_106_2_groupi_n_346 ^ csa_tree_add_106_2_groupi_n_345);
 assign csa_tree_add_106_2_groupi_n_633 = ~(csa_tree_add_106_2_groupi_n_434 & csa_tree_add_106_2_groupi_n_632);
 assign csa_tree_add_106_2_groupi_n_630 = (csa_tree_add_106_2_groupi_n_332 & csa_tree_add_106_2_groupi_n_333);
 assign csa_tree_add_106_2_groupi_n_631 = (csa_tree_add_106_2_groupi_n_332 ^ csa_tree_add_106_2_groupi_n_333);
 assign csa_tree_add_106_2_groupi_n_617 = ~(csa_tree_add_106_2_groupi_n_432 | csa_tree_add_106_2_groupi_n_44);
 assign csa_tree_add_106_2_groupi_n_605 = ~(csa_tree_add_106_2_groupi_n_428 | csa_tree_add_106_2_groupi_n_39);
 assign csa_tree_add_106_2_groupi_n_603 = ~((n_1499 | csa_tree_add_106_2_groupi_n_92) & (csa_tree_add_106_2_groupi_n_312
    | csa_tree_add_106_2_groupi_n_46));
 assign csa_tree_add_106_2_groupi_n_602 = ~((n_1499 | csa_tree_add_106_2_groupi_n_311) & (csa_tree_add_106_2_groupi_n_240
    | csa_tree_add_106_2_groupi_n_46));
 assign csa_tree_add_106_2_groupi_n_599 = ~((n_1499 | csa_tree_add_106_2_groupi_n_240) & (csa_tree_add_106_2_groupi_n_248
    | csa_tree_add_106_2_groupi_n_46));
 assign csa_tree_add_106_2_groupi_n_592 = ~((n_1499 | csa_tree_add_106_2_groupi_n_312) & (csa_tree_add_106_2_groupi_n_311
    | csa_tree_add_106_2_groupi_n_46));
 assign csa_tree_add_106_2_groupi_n_584 = ~(csa_tree_add_106_2_groupi_n_433 | csa_tree_add_106_2_groupi_n_43);
 assign csa_tree_add_106_2_groupi_n_563 = ~((csa_tree_add_106_2_groupi_n_343 | csa_tree_add_106_2_groupi_n_131)
    & (csa_tree_add_106_2_groupi_n_226 | csa_tree_add_106_2_groupi_n_126));
 assign csa_tree_add_106_2_groupi_n_558 = ~((csa_tree_add_106_2_groupi_n_343 | csa_tree_add_106_2_groupi_n_126)
    & (csa_tree_add_106_2_groupi_n_226 | csa_tree_add_106_2_groupi_n_119));
 assign csa_tree_add_106_2_groupi_n_554 = ~((csa_tree_add_106_2_groupi_n_344 | csa_tree_add_106_2_groupi_n_86)
    & (csa_tree_add_106_2_groupi_n_225 | csa_tree_add_106_2_groupi_n_113));
 assign csa_tree_add_106_2_groupi_n_553 = ~((csa_tree_add_106_2_groupi_n_343 | csa_tree_add_106_2_groupi_n_87)
    & (csa_tree_add_106_2_groupi_n_226 | csa_tree_add_106_2_groupi_n_131));
 assign csa_tree_add_106_2_groupi_n_538 = ~(csa_tree_add_106_2_groupi_n_429 | csa_tree_add_106_2_groupi_n_41);
 assign csa_tree_add_106_2_groupi_n_536 = ~(csa_tree_add_106_2_groupi_n_430 | csa_tree_add_106_2_groupi_n_7);
 assign csa_tree_add_106_2_groupi_n_534 = ~(csa_tree_add_106_2_groupi_n_431 | csa_tree_add_106_2_groupi_n_42);
 assign csa_tree_add_106_2_groupi_n_504 = ~((csa_tree_add_106_2_groupi_n_1 | csa_tree_add_106_2_groupi_n_153)
    & (csa_tree_add_106_2_groupi_n_224 | csa_tree_add_106_2_groupi_n_170));
 assign csa_tree_add_106_2_groupi_n_503 = ~((csa_tree_add_106_2_groupi_n_1 | csa_tree_add_106_2_groupi_n_161)
    & (csa_tree_add_106_2_groupi_n_224 | csa_tree_add_106_2_groupi_n_153));
 assign csa_tree_add_106_2_groupi_n_497 = ~((csa_tree_add_106_2_groupi_n_2 | csa_tree_add_106_2_groupi_n_187)
    & (csa_tree_add_106_2_groupi_n_223 | csa_tree_add_106_2_groupi_n_177));
 assign csa_tree_add_106_2_groupi_n_496 = ~((csa_tree_add_106_2_groupi_n_2 | csa_tree_add_106_2_groupi_n_89)
    & (csa_tree_add_106_2_groupi_n_223 | csa_tree_add_106_2_groupi_n_187));
 assign csa_tree_add_106_2_groupi_n_491 = ~((csa_tree_add_106_2_groupi_n_1 | csa_tree_add_106_2_groupi_n_88)
    & (csa_tree_add_106_2_groupi_n_224 | csa_tree_add_106_2_groupi_n_161));
 assign csa_tree_add_106_2_groupi_n_465 = ~((csa_tree_add_106_2_groupi_n_4 | csa_tree_add_106_2_groupi_n_203)
    & (csa_tree_add_106_2_groupi_n_221 | csa_tree_add_106_2_groupi_n_94));
 assign csa_tree_add_106_2_groupi_n_463 = ~((csa_tree_add_106_2_groupi_n_4 | csa_tree_add_106_2_groupi_n_90)
    & (csa_tree_add_106_2_groupi_n_221 | csa_tree_add_106_2_groupi_n_195));
 assign csa_tree_add_106_2_groupi_n_462 = ~((csa_tree_add_106_2_groupi_n_4 | csa_tree_add_106_2_groupi_n_195)
    & (csa_tree_add_106_2_groupi_n_221 | csa_tree_add_106_2_groupi_n_203));
 assign csa_tree_add_106_2_groupi_n_455 = ~((csa_tree_add_106_2_groupi_n_3 | csa_tree_add_106_2_groupi_n_91)
    & (csa_tree_add_106_2_groupi_n_222 | csa_tree_add_106_2_groupi_n_245));
 assign csa_tree_add_106_2_groupi_n_437 = ~((csa_tree_add_106_2_groupi_n_3 | csa_tree_add_106_2_groupi_n_245)
    & (csa_tree_add_106_2_groupi_n_222 | csa_tree_add_106_2_groupi_n_233));
 assign csa_tree_add_106_2_groupi_n_433 = ~((csa_tree_add_106_2_groupi_n_79 & csa_tree_add_106_2_groupi_n_47)
    | (csa_tree_add_106_2_groupi_n_42 & csa_tree_add_106_2_groupi_n_34));
 assign csa_tree_add_106_2_groupi_n_432 = ~((csa_tree_add_106_2_groupi_n_78 & csa_tree_add_106_2_groupi_n_8)
    | (csa_tree_add_106_2_groupi_n_7 & csa_tree_add_106_2_groupi_n_37));
 assign csa_tree_add_106_2_groupi_n_431 = ~((csa_tree_add_106_2_groupi_n_80 & csa_tree_add_106_2_groupi_n_47)
    | (csa_tree_add_106_2_groupi_n_41 & csa_tree_add_106_2_groupi_n_35));
 assign csa_tree_add_106_2_groupi_n_430 = ~((csa_tree_add_106_2_groupi_n_82 & csa_tree_add_106_2_groupi_n_8)
    | (csa_tree_add_106_2_groupi_n_39 & csa_tree_add_106_2_groupi_n_74));
 assign csa_tree_add_106_2_groupi_n_429 = ~((csa_tree_add_106_2_groupi_n_81 & csa_tree_add_106_2_groupi_n_47)
    | (csa_tree_add_106_2_groupi_n_40 & csa_tree_add_106_2_groupi_n_73));
 assign csa_tree_add_106_2_groupi_n_428 = ~((csa_tree_add_106_2_groupi_n_83 & csa_tree_add_106_2_groupi_n_8)
    | (csa_tree_add_106_2_groupi_n_38 & csa_tree_add_106_2_groupi_n_36));
 assign csa_tree_add_106_2_groupi_n_427 = ~((csa_tree_add_106_2_groupi_n_335 & n_1413) | (csa_tree_add_106_2_groupi_n_229
    & n_1412));
 assign csa_tree_add_106_2_groupi_n_426 = ~((csa_tree_add_106_2_groupi_n_337 & n_1329) | (csa_tree_add_106_2_groupi_n_227
    & n_1328));
 assign csa_tree_add_106_2_groupi_n_434 = ~((csa_tree_add_106_2_groupi_n_337 & n_1330) | (csa_tree_add_106_2_groupi_n_227
    & n_1329));
 assign csa_tree_add_106_2_groupi_n_385 = ~((csa_tree_add_106_2_groupi_n_336 | csa_tree_add_106_2_groupi_n_8)
    & (csa_tree_add_106_2_groupi_n_230 | csa_tree_add_106_2_groupi_n_61));
 assign csa_tree_add_106_2_groupi_n_384 = ~((csa_tree_add_106_2_groupi_n_338 | csa_tree_add_106_2_groupi_n_47)
    & (csa_tree_add_106_2_groupi_n_228 | csa_tree_add_106_2_groupi_n_15));
 assign csa_tree_add_106_2_groupi_n_370 = ~((n_1492 | csa_tree_add_106_2_groupi_n_268) & (csa_tree_add_106_2_groupi_n_262
    | csa_tree_add_106_2_groupi_n_45));
 assign csa_tree_add_106_2_groupi_n_362 = ~((n_1492 | csa_tree_add_106_2_groupi_n_93) & (csa_tree_add_106_2_groupi_n_268
    | csa_tree_add_106_2_groupi_n_45));
 assign csa_tree_add_106_2_groupi_n_350 = ~(csa_tree_add_106_2_groupi_n_225 | csa_tree_add_106_2_groupi_n_8);
 assign csa_tree_add_106_2_groupi_n_349 = ~(csa_tree_add_106_2_groupi_n_226 | csa_tree_add_106_2_groupi_n_47);
 assign csa_tree_add_106_2_groupi_n_348 = ~(csa_tree_add_106_2_groupi_n_223 | csa_tree_add_106_2_groupi_n_8);
 assign csa_tree_add_106_2_groupi_n_347 = ~(csa_tree_add_106_2_groupi_n_224 | csa_tree_add_106_2_groupi_n_47);
 assign csa_tree_add_106_2_groupi_n_346 = ~(csa_tree_add_106_2_groupi_n_221 | csa_tree_add_106_2_groupi_n_47);
 assign csa_tree_add_106_2_groupi_n_345 = ~(csa_tree_add_106_2_groupi_n_222 | csa_tree_add_106_2_groupi_n_8);
 assign csa_tree_add_106_2_groupi_n_333 = ~(csa_tree_add_106_2_groupi_n_230 | csa_tree_add_106_2_groupi_n_8);
 assign csa_tree_add_106_2_groupi_n_332 = ~(csa_tree_add_106_2_groupi_n_228 | csa_tree_add_106_2_groupi_n_47);
 assign csa_tree_add_106_2_groupi_n_220 = ~((csa_tree_add_106_2_groupi_n_35 & n_1442) | (csa_tree_add_106_2_groupi_n_42
    & n_1443));
 assign csa_tree_add_106_2_groupi_n_218 = ~((csa_tree_add_106_2_groupi_n_36 & n_1435) | (csa_tree_add_106_2_groupi_n_39
    & n_1436));
 assign csa_tree_add_106_2_groupi_n_217 = ~((csa_tree_add_106_2_groupi_n_73 & n_1444) | (csa_tree_add_106_2_groupi_n_41
    & n_1445));
 assign csa_tree_add_106_2_groupi_n_215 = ~((csa_tree_add_106_2_groupi_n_74 & n_1433) | (csa_tree_add_106_2_groupi_n_7
    & n_1434));
 assign csa_tree_add_106_2_groupi_n_212 = ~((csa_tree_add_106_2_groupi_n_34 & n_1440) | (csa_tree_add_106_2_groupi_n_43
    & n_1441));
 assign csa_tree_add_106_2_groupi_n_211 = ~((csa_tree_add_106_2_groupi_n_37 & n_1431) | (csa_tree_add_106_2_groupi_n_44
    & n_1432));
 assign csa_tree_add_106_2_groupi_n_312 = ~((csa_tree_add_106_2_groupi_n_40 & n_1349) | (csa_tree_add_106_2_groupi_n_15
    & n_1446));
 assign csa_tree_add_106_2_groupi_n_311 = ~((csa_tree_add_106_2_groupi_n_40 & n_1348) | (csa_tree_add_106_2_groupi_n_21
    & n_1446));
 assign csa_tree_add_106_2_groupi_n_268 = ~((csa_tree_add_106_2_groupi_n_38 & n_1428) | (csa_tree_add_106_2_groupi_n_61
    & n_1437));
 assign csa_tree_add_106_2_groupi_n_245 = ~((csa_tree_add_106_2_groupi_n_39 & n_1428) | (csa_tree_add_106_2_groupi_n_61
    & n_1435));
 assign csa_tree_add_106_2_groupi_n_240 = ~((csa_tree_add_106_2_groupi_n_40 & n_1347) | (csa_tree_add_106_2_groupi_n_48
    & n_1446));
 assign csa_tree_add_106_2_groupi_n_208 = ~(csa_tree_add_106_2_groupi_n_77 | csa_tree_add_106_2_groupi_n_40);
 assign csa_tree_add_106_2_groupi_n_207 = ~(csa_tree_add_106_2_groupi_n_76 | csa_tree_add_106_2_groupi_n_38);
 assign csa_tree_add_106_2_groupi_n_93 = ~((csa_tree_add_106_2_groupi_n_38 & n_1429) | (csa_tree_add_106_2_groupi_n_8
    & n_1437));
 assign csa_tree_add_106_2_groupi_n_92 = ~((csa_tree_add_106_2_groupi_n_40 & n_1350) | (csa_tree_add_106_2_groupi_n_47
    & n_1446));
 assign csa_tree_add_106_2_groupi_n_91 = ~((csa_tree_add_106_2_groupi_n_39 & n_1429) | (csa_tree_add_106_2_groupi_n_8
    & n_1435));
 assign csa_tree_add_106_2_groupi_n_90 = ~((csa_tree_add_106_2_groupi_n_41 & n_1350) | (csa_tree_add_106_2_groupi_n_47
    & n_1444));
 assign csa_tree_add_106_2_groupi_n_89 = ~((csa_tree_add_106_2_groupi_n_7 & n_1429) | (csa_tree_add_106_2_groupi_n_8
    & n_1433));
 assign csa_tree_add_106_2_groupi_n_88 = ~((csa_tree_add_106_2_groupi_n_42 & n_1350) | (csa_tree_add_106_2_groupi_n_47
    & n_1442));
 assign csa_tree_add_106_2_groupi_n_87 = ~((csa_tree_add_106_2_groupi_n_43 & n_1350) | (csa_tree_add_106_2_groupi_n_47
    & n_1440));
 assign csa_tree_add_106_2_groupi_n_86 = ~((csa_tree_add_106_2_groupi_n_44 & n_1429) | (csa_tree_add_106_2_groupi_n_8
    & n_1431));
 assign csa_tree_add_106_2_groupi_n_203 = ~((csa_tree_add_106_2_groupi_n_41 & n_1348) | (csa_tree_add_106_2_groupi_n_21
    & n_1444));
 assign csa_tree_add_106_2_groupi_n_195 = ~((csa_tree_add_106_2_groupi_n_41 & n_1349) | (csa_tree_add_106_2_groupi_n_15
    & n_1444));
 assign csa_tree_add_106_2_groupi_n_187 = ~((csa_tree_add_106_2_groupi_n_7 & n_1428) | (csa_tree_add_106_2_groupi_n_61
    & n_1433));
 assign csa_tree_add_106_2_groupi_n_161 = ~((csa_tree_add_106_2_groupi_n_42 & n_1349) | (csa_tree_add_106_2_groupi_n_15
    & n_1442));
 assign csa_tree_add_106_2_groupi_n_153 = ~((csa_tree_add_106_2_groupi_n_42 & n_1348) | (csa_tree_add_106_2_groupi_n_21
    & n_1442));
 assign csa_tree_add_106_2_groupi_n_131 = ~((csa_tree_add_106_2_groupi_n_43 & n_1349) | (csa_tree_add_106_2_groupi_n_15
    & n_1440));
 assign csa_tree_add_106_2_groupi_n_126 = ~((csa_tree_add_106_2_groupi_n_43 & n_1348) | (csa_tree_add_106_2_groupi_n_21
    & n_1440));
 assign csa_tree_add_106_2_groupi_n_83 = ~(n_1437 & n_1436);
 assign csa_tree_add_106_2_groupi_n_82 = ~(n_1435 & n_1434);
 assign csa_tree_add_106_2_groupi_n_81 = ~(n_1446 & n_1445);
 assign csa_tree_add_106_2_groupi_n_80 = ~(n_1444 & n_1443);
 assign csa_tree_add_106_2_groupi_n_79 = ~(n_1442 & n_1441);
 assign csa_tree_add_106_2_groupi_n_78 = ~(n_1433 & n_1432);
 assign csa_tree_add_106_2_groupi_n_77 = ~(csa_tree_add_106_2_groupi_n_46 | csa_tree_add_106_2_groupi_n_47);
 assign csa_tree_add_106_2_groupi_n_76 = ~(csa_tree_add_106_2_groupi_n_45 | csa_tree_add_106_2_groupi_n_8);
 assign csa_tree_add_106_2_groupi_n_74 = ~n_1434;
 assign csa_tree_add_106_2_groupi_n_73 = ~n_1445;
 assign csa_tree_add_106_2_groupi_n_72 = ~n_1411;
 assign csa_tree_add_106_2_groupi_n_71 = ~n_1326;
 assign csa_tree_add_106_2_groupi_n_70 = ~n_1327;
 assign csa_tree_add_106_2_groupi_n_69 = ~n_1412;
 assign csa_tree_add_106_2_groupi_n_68 = ~n_1413;
 assign csa_tree_add_106_2_groupi_n_65 = ~n_1425;
 assign csa_tree_add_106_2_groupi_n_64 = ~n_1422;
 assign csa_tree_add_106_2_groupi_n_62 = ~n_1424;
 assign csa_tree_add_106_2_groupi_n_61 = ~n_1428;
 assign csa_tree_add_106_2_groupi_n_58 = ~n_1331;
 assign csa_tree_add_106_2_groupi_n_53 = ~n_1427;
 assign csa_tree_add_106_2_groupi_n_52 = ~n_1333;
 assign csa_tree_add_106_2_groupi_n_51 = ~n_1423;
 assign csa_tree_add_106_2_groupi_n_49 = ~n_1426;
 assign csa_tree_add_106_2_groupi_n_47 = ~n_1350;
 assign csa_tree_add_106_2_groupi_n_37 = ~n_1432;
 assign csa_tree_add_106_2_groupi_n_36 = ~n_1436;
 assign csa_tree_add_106_2_groupi_n_35 = ~n_1443;
 assign csa_tree_add_106_2_groupi_n_34 = ~n_1441;
 assign csa_tree_add_106_2_groupi_n_32 = ~n_1328;
 assign csa_tree_add_106_2_groupi_n_31 = ~n_1332;
 assign csa_tree_add_106_2_groupi_n_24 = ~n_1335;
 assign csa_tree_add_106_2_groupi_n_23 = ~n_1329;
 assign csa_tree_add_106_2_groupi_n_22 = ~n_1421;
 assign csa_tree_add_106_2_groupi_n_20 = ~n_1334;
 assign csa_tree_add_106_2_groupi_n_19 = ~n_1330;
 assign csa_tree_add_106_2_groupi_n_17 = ~n_1418;
 assign csa_tree_add_106_2_groupi_n_16 = ~n_1414;
 assign csa_tree_add_106_2_groupi_n_14 = ~n_1415;
 assign csa_tree_add_106_2_groupi_n_13 = ~n_1416;
 assign csa_tree_add_106_2_groupi_n_12 = ~n_1420;
 assign csa_tree_add_106_2_groupi_n_11 = ~n_1417;
 assign csa_tree_add_106_2_groupi_n_9 = ~n_1419;
 assign csa_tree_add_106_2_groupi_n_8 = ~n_1429;
 assign csa_tree_mul_77_11_groupi_n_11 = ~(csa_tree_mul_77_11_groupi_n_563 | ~csa_tree_mul_77_11_groupi_n_552);
 assign n_1324 = ~(csa_tree_mul_77_11_groupi_n_619 ^ csa_tree_mul_77_11_groupi_n_386);
 assign n_1325 = ~(csa_tree_mul_77_11_groupi_n_621 ^ csa_tree_mul_77_11_groupi_n_419);
 assign n_1326 = ~(csa_tree_mul_77_11_groupi_n_620 ^ csa_tree_mul_77_11_groupi_n_448);
 assign n_1328 = ~(csa_tree_mul_77_11_groupi_n_609 ^ csa_tree_mul_77_11_groupi_n_515);
 assign n_1329 = ~(csa_tree_mul_77_11_groupi_n_615 ^ csa_tree_mul_77_11_groupi_n_506);
 assign n_1330 = ~(csa_tree_mul_77_11_groupi_n_614 ^ csa_tree_mul_77_11_groupi_n_512);
 assign n_1332 = ~(csa_tree_mul_77_11_groupi_n_613 ^ csa_tree_mul_77_11_groupi_n_510);
 assign csa_tree_mul_77_11_groupi_n_621 = ~(csa_tree_mul_77_11_groupi_n_514 | (csa_tree_mul_77_11_groupi_n_608
    & csa_tree_mul_77_11_groupi_n_487));
 assign csa_tree_mul_77_11_groupi_n_620 = ~(csa_tree_mul_77_11_groupi_n_460 & (csa_tree_mul_77_11_groupi_n_607
    | csa_tree_mul_77_11_groupi_n_459));
 assign n_1327 = ~(csa_tree_mul_77_11_groupi_n_607 ^ csa_tree_mul_77_11_groupi_n_481);
 assign csa_tree_mul_77_11_groupi_n_617 = ~(csa_tree_mul_77_11_groupi_n_601 | (csa_tree_mul_77_11_groupi_n_606
    & csa_tree_mul_77_11_groupi_n_522));
 assign csa_tree_mul_77_11_groupi_n_615 = ~(csa_tree_mul_77_11_groupi_n_533 | (csa_tree_mul_77_11_groupi_n_605
    & csa_tree_mul_77_11_groupi_n_518));
 assign csa_tree_mul_77_11_groupi_n_614 = ~(csa_tree_mul_77_11_groupi_n_495 & ~(csa_tree_mul_77_11_groupi_n_605
    & csa_tree_mul_77_11_groupi_n_498));
 assign n_1331 = ~(csa_tree_mul_77_11_groupi_n_605 ^ csa_tree_mul_77_11_groupi_n_511);
 assign n_1333 = ~(csa_tree_mul_77_11_groupi_n_604 ^ csa_tree_mul_77_11_groupi_n_509);
 assign n_1334 = ~(csa_tree_mul_77_11_groupi_n_603 ^ csa_tree_mul_77_11_groupi_n_554);
 assign csa_tree_mul_77_11_groupi_n_609 = ~(csa_tree_mul_77_11_groupi_n_497 & (csa_tree_mul_77_11_groupi_n_585
    & (csa_tree_mul_77_11_groupi_n_536 | csa_tree_mul_77_11_groupi_n_600)));
 assign csa_tree_mul_77_11_groupi_n_608 = ~csa_tree_mul_77_11_groupi_n_607;
 assign csa_tree_mul_77_11_groupi_n_607 = ~(csa_tree_mul_77_11_groupi_n_606 | csa_tree_mul_77_11_groupi_n_590);
 assign csa_tree_mul_77_11_groupi_n_606 = ~(csa_tree_mul_77_11_groupi_n_544 | csa_tree_mul_77_11_groupi_n_600);
 assign csa_tree_mul_77_11_groupi_n_605 = ~(csa_tree_mul_77_11_groupi_n_600 & ~csa_tree_mul_77_11_groupi_n_575);
 assign n_1335 = ~(csa_tree_mul_77_11_groupi_n_594 ^ csa_tree_mul_77_11_groupi_n_553);
 assign csa_tree_mul_77_11_groupi_n_593 = ~(csa_tree_mul_77_11_groupi_n_531 | (csa_tree_mul_77_11_groupi_n_583
    & csa_tree_mul_77_11_groupi_n_513));
 assign csa_tree_mul_77_11_groupi_n_592 = ~(csa_tree_mul_77_11_groupi_n_483 & ~(csa_tree_mul_77_11_groupi_n_583
    & csa_tree_mul_77_11_groupi_n_485));
 assign csa_tree_mul_77_11_groupi_n_591 = ~(csa_tree_mul_77_11_groupi_n_586 | ((csa_tree_mul_77_11_groupi_n_542
    & csa_tree_mul_77_11_groupi_n_539) | (csa_tree_mul_77_11_groupi_n_531 & csa_tree_mul_77_11_groupi_n_557)));
 assign csa_tree_mul_77_11_groupi_n_590 = ~(csa_tree_mul_77_11_groupi_n_488 & (csa_tree_mul_77_11_groupi_n_559
    & (csa_tree_mul_77_11_groupi_n_576 | csa_tree_mul_77_11_groupi_n_544)));
 assign csa_tree_mul_77_11_groupi_n_587 = ~(csa_tree_mul_77_11_groupi_n_538 & (csa_tree_mul_77_11_groupi_n_584
    & (csa_tree_mul_77_11_groupi_n_573 | csa_tree_mul_77_11_groupi_n_548)));
 assign csa_tree_mul_77_11_groupi_n_586 = ~(csa_tree_mul_77_11_groupi_n_534 & ~(csa_tree_mul_77_11_groupi_n_574
    & csa_tree_mul_77_11_groupi_n_565));
 assign csa_tree_mul_77_11_groupi_n_585 = ~((csa_tree_mul_77_11_groupi_n_518 & (csa_tree_mul_77_11_groupi_n_494
    & csa_tree_mul_77_11_groupi_n_575)) | (csa_tree_mul_77_11_groupi_n_533 & csa_tree_mul_77_11_groupi_n_494));
 assign csa_tree_mul_77_11_groupi_n_584 = ~((csa_tree_mul_77_11_groupi_n_513 & (csa_tree_mul_77_11_groupi_n_530
    & csa_tree_mul_77_11_groupi_n_574)) | (csa_tree_mul_77_11_groupi_n_531 & csa_tree_mul_77_11_groupi_n_530));
 assign csa_tree_mul_77_11_groupi_n_583 = ~csa_tree_mul_77_11_groupi_n_582;
 assign csa_tree_mul_77_11_groupi_n_582 = ~(csa_tree_mul_77_11_groupi_n_574 | ~csa_tree_mul_77_11_groupi_n_573);
 assign csa_tree_mul_77_11_groupi_n_581 = ~(csa_tree_mul_77_11_groupi_n_551 & (csa_tree_mul_77_11_groupi_n_571
    | csa_tree_mul_77_11_groupi_n_556));
 assign csa_tree_mul_77_11_groupi_n_576 = ~csa_tree_mul_77_11_groupi_n_575;
 assign csa_tree_mul_77_11_groupi_n_574 = ~(csa_tree_mul_77_11_groupi_n_11 & ~(csa_tree_mul_77_11_groupi_n_568
    & csa_tree_mul_77_11_groupi_n_535));
 assign csa_tree_mul_77_11_groupi_n_573 = ~(csa_tree_mul_77_11_groupi_n_561 & csa_tree_mul_77_11_groupi_n_568);
 assign csa_tree_mul_77_11_groupi_n_572 = ~(csa_tree_mul_77_11_groupi_n_560 & csa_tree_mul_77_11_groupi_n_521);
 assign csa_tree_mul_77_11_groupi_n_571 = ~(csa_tree_mul_77_11_groupi_n_561 | csa_tree_mul_77_11_groupi_n_535);
 assign csa_tree_mul_77_11_groupi_n_570 = ~(csa_tree_mul_77_11_groupi_n_461 & (csa_tree_mul_77_11_groupi_n_549
    | csa_tree_mul_77_11_groupi_n_462));
 assign csa_tree_mul_77_11_groupi_n_568 = ~(csa_tree_mul_77_11_groupi_n_556 | csa_tree_mul_77_11_groupi_n_550);
 assign csa_tree_mul_77_11_groupi_n_567 = ~(csa_tree_mul_77_11_groupi_n_550 | ~csa_tree_mul_77_11_groupi_n_552);
 assign csa_tree_mul_77_11_groupi_n_566 = ~(csa_tree_mul_77_11_groupi_n_556 | ~csa_tree_mul_77_11_groupi_n_551);
 assign csa_tree_mul_77_11_groupi_n_565 = ~csa_tree_mul_77_11_groupi_n_564;
 assign csa_tree_mul_77_11_groupi_n_564 = ~(csa_tree_mul_77_11_groupi_n_557 & csa_tree_mul_77_11_groupi_n_513);
 assign csa_tree_mul_77_11_groupi_n_563 = ~(csa_tree_mul_77_11_groupi_n_551 | csa_tree_mul_77_11_groupi_n_550);
 assign csa_tree_mul_77_11_groupi_n_561 = ~(csa_tree_mul_77_11_groupi_n_500 | (csa_tree_mul_77_11_groupi_n_462
    | csa_tree_mul_77_11_groupi_n_549));
 assign csa_tree_mul_77_11_groupi_n_559 = ~(csa_tree_mul_77_11_groupi_n_517 | (csa_tree_mul_77_11_groupi_n_533
    & csa_tree_mul_77_11_groupi_n_520));
 assign csa_tree_mul_77_11_groupi_n_555 = ~(csa_tree_mul_77_11_groupi_n_542 & csa_tree_mul_77_11_groupi_n_534);
 assign csa_tree_mul_77_11_groupi_n_557 = (csa_tree_mul_77_11_groupi_n_542 & csa_tree_mul_77_11_groupi_n_530);
 assign csa_tree_mul_77_11_groupi_n_556 = ~(csa_tree_mul_77_11_groupi_n_546 | csa_tree_mul_77_11_groupi_n_477);
 assign csa_tree_mul_77_11_groupi_n_548 = ~(csa_tree_mul_77_11_groupi_n_513 & csa_tree_mul_77_11_groupi_n_530);
 assign csa_tree_mul_77_11_groupi_n_547 = ~(csa_tree_mul_77_11_groupi_n_539 | ~csa_tree_mul_77_11_groupi_n_530);
 assign csa_tree_mul_77_11_groupi_n_552 = ~(csa_tree_mul_77_11_groupi_n_480 & csa_tree_mul_77_11_groupi_n_545);
 assign csa_tree_mul_77_11_groupi_n_551 = ~(csa_tree_mul_77_11_groupi_n_546 & csa_tree_mul_77_11_groupi_n_477);
 assign csa_tree_mul_77_11_groupi_n_550 = ~(csa_tree_mul_77_11_groupi_n_480 | csa_tree_mul_77_11_groupi_n_545);
 assign csa_tree_mul_77_11_groupi_n_549 = ~(csa_tree_mul_77_11_groupi_n_528 | csa_tree_mul_77_11_groupi_n_527);
 assign csa_tree_mul_77_11_groupi_n_538 = ~csa_tree_mul_77_11_groupi_n_539;
 assign csa_tree_mul_77_11_groupi_n_545 = ((csa_tree_mul_77_11_groupi_n_414 & csa_tree_mul_77_11_groupi_n_338)
    | ((csa_tree_mul_77_11_groupi_n_338 & csa_tree_mul_77_11_groupi_n_438) | (csa_tree_mul_77_11_groupi_n_438
    & csa_tree_mul_77_11_groupi_n_414)));
 assign csa_tree_mul_77_11_groupi_n_546 = (csa_tree_mul_77_11_groupi_n_338 ^ (csa_tree_mul_77_11_groupi_n_438
    ^ csa_tree_mul_77_11_groupi_n_414));
 assign csa_tree_mul_77_11_groupi_n_537 = ~(csa_tree_mul_77_11_groupi_n_514 & csa_tree_mul_77_11_groupi_n_428);
 assign csa_tree_mul_77_11_groupi_n_544 = ~(csa_tree_mul_77_11_groupi_n_518 & csa_tree_mul_77_11_groupi_n_520);
 assign csa_tree_mul_77_11_groupi_n_536 = ~(csa_tree_mul_77_11_groupi_n_518 & csa_tree_mul_77_11_groupi_n_494);
 assign csa_tree_mul_77_11_groupi_n_542 = (csa_tree_mul_77_11_groupi_n_505 | csa_tree_mul_77_11_groupi_n_523);
 assign csa_tree_mul_77_11_groupi_n_539 = (csa_tree_mul_77_11_groupi_n_524 & csa_tree_mul_77_11_groupi_n_471);
 assign csa_tree_mul_77_11_groupi_n_528 = ~(csa_tree_mul_77_11_groupi_n_493 & (csa_tree_mul_77_11_groupi_n_5
    | csa_tree_mul_77_11_groupi_n_430));
 assign csa_tree_mul_77_11_groupi_n_527 = ~(csa_tree_mul_77_11_groupi_n_464 & (csa_tree_mul_77_11_groupi_n_5
    | csa_tree_mul_77_11_groupi_n_418));
 assign csa_tree_mul_77_11_groupi_n_535 = ~(csa_tree_mul_77_11_groupi_n_490 & (csa_tree_mul_77_11_groupi_n_500
    | csa_tree_mul_77_11_groupi_n_461));
 assign csa_tree_mul_77_11_groupi_n_534 = ~(csa_tree_mul_77_11_groupi_n_505 & csa_tree_mul_77_11_groupi_n_523);
 assign csa_tree_mul_77_11_groupi_n_533 = ~(csa_tree_mul_77_11_groupi_n_503 & (csa_tree_mul_77_11_groupi_n_495
    | csa_tree_mul_77_11_groupi_n_499));
 assign csa_tree_mul_77_11_groupi_n_531 = ~(csa_tree_mul_77_11_groupi_n_489 & (csa_tree_mul_77_11_groupi_n_484
    | csa_tree_mul_77_11_groupi_n_483));
 assign csa_tree_mul_77_11_groupi_n_530 = (csa_tree_mul_77_11_groupi_n_524 | csa_tree_mul_77_11_groupi_n_471);
 assign csa_tree_mul_77_11_groupi_n_525 = ((csa_tree_mul_77_11_groupi_n_427 & csa_tree_mul_77_11_groupi_n_361)
    | ((csa_tree_mul_77_11_groupi_n_361 & csa_tree_mul_77_11_groupi_n_422) | (csa_tree_mul_77_11_groupi_n_422
    & csa_tree_mul_77_11_groupi_n_427)));
 assign csa_tree_mul_77_11_groupi_n_526 = (csa_tree_mul_77_11_groupi_n_361 ^ (csa_tree_mul_77_11_groupi_n_422
    ^ csa_tree_mul_77_11_groupi_n_427));
 assign csa_tree_mul_77_11_groupi_n_523 = ((csa_tree_mul_77_11_groupi_n_425 & csa_tree_mul_77_11_groupi_n_420)
    | ((csa_tree_mul_77_11_groupi_n_420 & csa_tree_mul_77_11_groupi_n_374) | (csa_tree_mul_77_11_groupi_n_374
    & csa_tree_mul_77_11_groupi_n_425)));
 assign csa_tree_mul_77_11_groupi_n_524 = (csa_tree_mul_77_11_groupi_n_420 ^ (csa_tree_mul_77_11_groupi_n_374
    ^ csa_tree_mul_77_11_groupi_n_425));
 assign csa_tree_mul_77_11_groupi_n_517 = ~(csa_tree_mul_77_11_groupi_n_497 | csa_tree_mul_77_11_groupi_n_501);
 assign csa_tree_mul_77_11_groupi_n_522 = (csa_tree_mul_77_11_groupi_n_487 & csa_tree_mul_77_11_groupi_n_428);
 assign csa_tree_mul_77_11_groupi_n_520 = ~(csa_tree_mul_77_11_groupi_n_501 | ~csa_tree_mul_77_11_groupi_n_494);
 assign csa_tree_mul_77_11_groupi_n_515 = ~(csa_tree_mul_77_11_groupi_n_488 & ~csa_tree_mul_77_11_groupi_n_501);
 assign csa_tree_mul_77_11_groupi_n_518 = ~(csa_tree_mul_77_11_groupi_n_499 | ~csa_tree_mul_77_11_groupi_n_498);
 assign csa_tree_mul_77_11_groupi_n_512 = ~(csa_tree_mul_77_11_groupi_n_503 & ~csa_tree_mul_77_11_groupi_n_499);
 assign csa_tree_mul_77_11_groupi_n_511 = ~(csa_tree_mul_77_11_groupi_n_498 & csa_tree_mul_77_11_groupi_n_495);
 assign csa_tree_mul_77_11_groupi_n_508 = ~(csa_tree_mul_77_11_groupi_n_484 | ~csa_tree_mul_77_11_groupi_n_489);
 assign csa_tree_mul_77_11_groupi_n_507 = ~(csa_tree_mul_77_11_groupi_n_486 | ~csa_tree_mul_77_11_groupi_n_483);
 assign csa_tree_mul_77_11_groupi_n_506 = (csa_tree_mul_77_11_groupi_n_494 & csa_tree_mul_77_11_groupi_n_497);
 assign csa_tree_mul_77_11_groupi_n_513 = ~(csa_tree_mul_77_11_groupi_n_484 | csa_tree_mul_77_11_groupi_n_486);
 assign csa_tree_mul_77_11_groupi_n_504 = ((csa_tree_mul_77_11_groupi_n_424 & csa_tree_mul_77_11_groupi_n_423)
    | ((csa_tree_mul_77_11_groupi_n_423 & csa_tree_mul_77_11_groupi_n_372) | (csa_tree_mul_77_11_groupi_n_372
    & csa_tree_mul_77_11_groupi_n_424)));
 assign csa_tree_mul_77_11_groupi_n_505 = (csa_tree_mul_77_11_groupi_n_423 ^ (csa_tree_mul_77_11_groupi_n_372
    ^ csa_tree_mul_77_11_groupi_n_424));
 assign csa_tree_mul_77_11_groupi_n_493 = ~(csa_tree_mul_77_11_groupi_n_3 & ~csa_tree_mul_77_11_groupi_n_440);
 assign csa_tree_mul_77_11_groupi_n_501 = ~(csa_tree_mul_77_11_groupi_n_457 | csa_tree_mul_77_11_groupi_n_473);
 assign csa_tree_mul_77_11_groupi_n_500 = ~(csa_tree_mul_77_11_groupi_n_478 | csa_tree_mul_77_11_groupi_n_454);
 assign csa_tree_mul_77_11_groupi_n_497 = ~(csa_tree_mul_77_11_groupi_n_474 & csa_tree_mul_77_11_groupi_n_469);
 assign csa_tree_mul_77_11_groupi_n_494 = (csa_tree_mul_77_11_groupi_n_474 | csa_tree_mul_77_11_groupi_n_469);
 assign csa_tree_mul_77_11_groupi_n_490 = ~csa_tree_mul_77_11_groupi_n_7;
 assign csa_tree_mul_77_11_groupi_n_485 = ~csa_tree_mul_77_11_groupi_n_486;
 assign csa_tree_mul_77_11_groupi_n_492 = ~(csa_tree_mul_77_11_groupi_n_3 & ~csa_tree_mul_77_11_groupi_n_463);
 assign csa_tree_mul_77_11_groupi_n_481 = ~(csa_tree_mul_77_11_groupi_n_459 | ~csa_tree_mul_77_11_groupi_n_460);
 assign csa_tree_mul_77_11_groupi_n_489 = ~(csa_tree_mul_77_11_groupi_n_472 & csa_tree_mul_77_11_groupi_n_449);
 assign csa_tree_mul_77_11_groupi_n_488 = ~(csa_tree_mul_77_11_groupi_n_457 & csa_tree_mul_77_11_groupi_n_473);
 assign csa_tree_mul_77_11_groupi_n_486 = ~(csa_tree_mul_77_11_groupi_n_450 | csa_tree_mul_77_11_groupi_n_479);
 assign csa_tree_mul_77_11_groupi_n_484 = ~(csa_tree_mul_77_11_groupi_n_472 | csa_tree_mul_77_11_groupi_n_449);
 assign csa_tree_mul_77_11_groupi_n_483 = ~(csa_tree_mul_77_11_groupi_n_450 & csa_tree_mul_77_11_groupi_n_479);
 assign csa_tree_mul_77_11_groupi_n_464 = ~csa_tree_mul_77_11_groupi_n_463;
 assign csa_tree_mul_77_11_groupi_n_479 = ((csa_tree_mul_77_11_groupi_n_413 & csa_tree_mul_77_11_groupi_n_381)
    | ((csa_tree_mul_77_11_groupi_n_381 & csa_tree_mul_77_11_groupi_n_363) | (csa_tree_mul_77_11_groupi_n_363
    & csa_tree_mul_77_11_groupi_n_413)));
 assign csa_tree_mul_77_11_groupi_n_480 = (csa_tree_mul_77_11_groupi_n_381 ^ (csa_tree_mul_77_11_groupi_n_363
    ^ csa_tree_mul_77_11_groupi_n_413));
 assign csa_tree_mul_77_11_groupi_n_477 = ((csa_tree_mul_77_11_groupi_n_439 & csa_tree_mul_77_11_groupi_n_277)
    | ((csa_tree_mul_77_11_groupi_n_277 & csa_tree_mul_77_11_groupi_n_403) | (csa_tree_mul_77_11_groupi_n_403
    & csa_tree_mul_77_11_groupi_n_439)));
 assign csa_tree_mul_77_11_groupi_n_478 = (csa_tree_mul_77_11_groupi_n_277 ^ (csa_tree_mul_77_11_groupi_n_403
    ^ csa_tree_mul_77_11_groupi_n_439));
 assign csa_tree_mul_77_11_groupi_n_475 = ((csa_tree_mul_77_11_groupi_n_426 & csa_tree_mul_77_11_groupi_n_350)
    | ((csa_tree_mul_77_11_groupi_n_350 & csa_tree_mul_77_11_groupi_n_398) | (csa_tree_mul_77_11_groupi_n_398
    & csa_tree_mul_77_11_groupi_n_426)));
 assign csa_tree_mul_77_11_groupi_n_476 = (csa_tree_mul_77_11_groupi_n_350 ^ (csa_tree_mul_77_11_groupi_n_398
    ^ csa_tree_mul_77_11_groupi_n_426));
 assign csa_tree_mul_77_11_groupi_n_471 = ((csa_tree_mul_77_11_groupi_n_421 & csa_tree_mul_77_11_groupi_n_388)
    | ((csa_tree_mul_77_11_groupi_n_388 & csa_tree_mul_77_11_groupi_n_379) | (csa_tree_mul_77_11_groupi_n_379
    & csa_tree_mul_77_11_groupi_n_421)));
 assign csa_tree_mul_77_11_groupi_n_472 = (csa_tree_mul_77_11_groupi_n_388 ^ (csa_tree_mul_77_11_groupi_n_379
    ^ csa_tree_mul_77_11_groupi_n_421));
 assign csa_tree_mul_77_11_groupi_n_463 = ~(csa_tree_mul_77_11_groupi_n_444 | ~csa_tree_mul_77_11_groupi_n_385);
 assign csa_tree_mul_77_11_groupi_n_462 = ~(csa_tree_mul_77_11_groupi_n_455 | csa_tree_mul_77_11_groupi_n_445);
 assign csa_tree_mul_77_11_groupi_n_461 = ~(csa_tree_mul_77_11_groupi_n_455 & csa_tree_mul_77_11_groupi_n_445);
 assign csa_tree_mul_77_11_groupi_n_454 = ((csa_tree_mul_77_11_groupi_n_404 & csa_tree_mul_77_11_groupi_n_255)
    | ((csa_tree_mul_77_11_groupi_n_255 & csa_tree_mul_77_11_groupi_n_377) | (csa_tree_mul_77_11_groupi_n_377
    & csa_tree_mul_77_11_groupi_n_404)));
 assign csa_tree_mul_77_11_groupi_n_455 = (csa_tree_mul_77_11_groupi_n_255 ^ (csa_tree_mul_77_11_groupi_n_377
    ^ csa_tree_mul_77_11_groupi_n_404));
 assign csa_tree_mul_77_11_groupi_n_452 = ((csa_tree_mul_77_11_groupi_n_396 & csa_tree_mul_77_11_groupi_n_355)
    | ((csa_tree_mul_77_11_groupi_n_355 & csa_tree_mul_77_11_groupi_n_397) | (csa_tree_mul_77_11_groupi_n_397
    & csa_tree_mul_77_11_groupi_n_396)));
 assign csa_tree_mul_77_11_groupi_n_453 = (csa_tree_mul_77_11_groupi_n_355 ^ (csa_tree_mul_77_11_groupi_n_397
    ^ csa_tree_mul_77_11_groupi_n_396));
 assign csa_tree_mul_77_11_groupi_n_451 = ~(csa_tree_mul_77_11_groupi_n_440 & (csa_tree_mul_77_11_groupi_n_441
    | csa_tree_mul_77_11_groupi_n_442));
 assign csa_tree_mul_77_11_groupi_n_449 = ((csa_tree_mul_77_11_groupi_n_380 & csa_tree_mul_77_11_groupi_n_389)
    | ((csa_tree_mul_77_11_groupi_n_389 & csa_tree_mul_77_11_groupi_n_353) | (csa_tree_mul_77_11_groupi_n_353
    & csa_tree_mul_77_11_groupi_n_380)));
 assign csa_tree_mul_77_11_groupi_n_450 = (csa_tree_mul_77_11_groupi_n_389 ^ (csa_tree_mul_77_11_groupi_n_353
    ^ csa_tree_mul_77_11_groupi_n_380));
 assign csa_tree_mul_77_11_groupi_n_447 = ~(csa_tree_mul_77_11_groupi_n_442 | ~csa_tree_mul_77_11_groupi_n_440);
 assign csa_tree_mul_77_11_groupi_n_445 = ~(csa_tree_mul_77_11_groupi_n_435 & ~(csa_tree_mul_77_11_groupi_n_365
    & csa_tree_mul_77_11_groupi_n_295));
 assign csa_tree_mul_77_11_groupi_n_444 = (csa_tree_mul_77_11_groupi_n_2 ^ csa_tree_mul_77_11_groupi_n_433);
 assign csa_tree_mul_77_11_groupi_n_438 = ((csa_tree_mul_77_11_groupi_n_339 & csa_tree_mul_77_11_groupi_n_206)
    | ((csa_tree_mul_77_11_groupi_n_206 & csa_tree_mul_77_11_groupi_n_358) | (csa_tree_mul_77_11_groupi_n_358
    & csa_tree_mul_77_11_groupi_n_339)));
 assign csa_tree_mul_77_11_groupi_n_439 = (csa_tree_mul_77_11_groupi_n_206 ^ (csa_tree_mul_77_11_groupi_n_358
    ^ csa_tree_mul_77_11_groupi_n_339));
 assign csa_tree_mul_77_11_groupi_n_442 = ~(csa_tree_mul_77_11_groupi_n_434 | csa_tree_mul_77_11_groupi_n_383);
 assign csa_tree_mul_77_11_groupi_n_441 = ~(csa_tree_mul_77_11_groupi_n_417 | csa_tree_mul_77_11_groupi_n_429);
 assign csa_tree_mul_77_11_groupi_n_440 = ~(csa_tree_mul_77_11_groupi_n_434 & csa_tree_mul_77_11_groupi_n_383);
 assign csa_tree_mul_77_11_groupi_n_435 = ~(csa_tree_mul_77_11_groupi_n_433 & (csa_tree_mul_77_11_groupi_n_365
    | csa_tree_mul_77_11_groupi_n_295));
 assign csa_tree_mul_77_11_groupi_n_430 = ~csa_tree_mul_77_11_groupi_n_429;
 assign csa_tree_mul_77_11_groupi_n_426 = ((csa_tree_mul_77_11_groupi_n_371 & csa_tree_mul_77_11_groupi_n_209)
    | ((csa_tree_mul_77_11_groupi_n_209 & csa_tree_mul_77_11_groupi_n_310) | (csa_tree_mul_77_11_groupi_n_310
    & csa_tree_mul_77_11_groupi_n_371)));
 assign csa_tree_mul_77_11_groupi_n_427 = (csa_tree_mul_77_11_groupi_n_209 ^ (csa_tree_mul_77_11_groupi_n_310
    ^ csa_tree_mul_77_11_groupi_n_371));
 assign csa_tree_mul_77_11_groupi_n_424 = ((csa_tree_mul_77_11_groupi_n_378 & csa_tree_mul_77_11_groupi_n_276)
    | ((csa_tree_mul_77_11_groupi_n_276 & csa_tree_mul_77_11_groupi_n_323) | (csa_tree_mul_77_11_groupi_n_323
    & csa_tree_mul_77_11_groupi_n_378)));
 assign csa_tree_mul_77_11_groupi_n_425 = (csa_tree_mul_77_11_groupi_n_276 ^ (csa_tree_mul_77_11_groupi_n_323
    ^ csa_tree_mul_77_11_groupi_n_378));
 assign csa_tree_mul_77_11_groupi_n_433 = ((csa_tree_mul_77_11_groupi_n_351 & csa_tree_mul_77_11_groupi_n_281)
    | ((csa_tree_mul_77_11_groupi_n_281 & csa_tree_mul_77_11_groupi_n_220) | (csa_tree_mul_77_11_groupi_n_220
    & csa_tree_mul_77_11_groupi_n_351)));
 assign csa_tree_mul_77_11_groupi_n_434 = (csa_tree_mul_77_11_groupi_n_281 ^ (csa_tree_mul_77_11_groupi_n_220
    ^ csa_tree_mul_77_11_groupi_n_351));
 assign csa_tree_mul_77_11_groupi_n_422 = ((csa_tree_mul_77_11_groupi_n_373 & csa_tree_mul_77_11_groupi_n_225)
    | ((csa_tree_mul_77_11_groupi_n_225 & csa_tree_mul_77_11_groupi_n_311) | (csa_tree_mul_77_11_groupi_n_311
    & csa_tree_mul_77_11_groupi_n_373)));
 assign csa_tree_mul_77_11_groupi_n_423 = (csa_tree_mul_77_11_groupi_n_225 ^ (csa_tree_mul_77_11_groupi_n_311
    ^ csa_tree_mul_77_11_groupi_n_373));
 assign csa_tree_mul_77_11_groupi_n_420 = ((csa_tree_mul_77_11_groupi_n_352 & csa_tree_mul_77_11_groupi_n_286)
    | ((csa_tree_mul_77_11_groupi_n_286 & csa_tree_mul_77_11_groupi_n_191) | (csa_tree_mul_77_11_groupi_n_191
    & csa_tree_mul_77_11_groupi_n_352)));
 assign csa_tree_mul_77_11_groupi_n_421 = (csa_tree_mul_77_11_groupi_n_286 ^ (csa_tree_mul_77_11_groupi_n_191
    ^ csa_tree_mul_77_11_groupi_n_352));
 assign csa_tree_mul_77_11_groupi_n_429 = ~(csa_tree_mul_77_11_groupi_n_387 | csa_tree_mul_77_11_groupi_n_412);
 assign csa_tree_mul_77_11_groupi_n_418 = ~csa_tree_mul_77_11_groupi_n_417;
 assign csa_tree_mul_77_11_groupi_n_417 = ~(csa_tree_mul_77_11_groupi_n_405 & (csa_tree_mul_77_11_groupi_n_387
    | csa_tree_mul_77_11_groupi_n_364));
 assign csa_tree_mul_77_11_groupi_n_416 = ~(csa_tree_mul_77_11_groupi_n_412 & csa_tree_mul_77_11_groupi_n_364);
 assign csa_tree_mul_77_11_groupi_n_413 = ((csa_tree_mul_77_11_groupi_n_343 & csa_tree_mul_77_11_groupi_n_279)
    | ((csa_tree_mul_77_11_groupi_n_279 & csa_tree_mul_77_11_groupi_n_208) | (csa_tree_mul_77_11_groupi_n_208
    & csa_tree_mul_77_11_groupi_n_343)));
 assign csa_tree_mul_77_11_groupi_n_414 = (csa_tree_mul_77_11_groupi_n_279 ^ (csa_tree_mul_77_11_groupi_n_208
    ^ csa_tree_mul_77_11_groupi_n_343));
 assign csa_tree_mul_77_11_groupi_n_412 = ~(csa_tree_mul_77_11_groupi_n_406 & csa_tree_mul_77_11_groupi_n_344);
 assign csa_tree_mul_77_11_groupi_n_409 = ~(csa_tree_mul_77_11_groupi_n_405 & ~csa_tree_mul_77_11_groupi_n_387);
 assign csa_tree_mul_77_11_groupi_n_407 = ((csa_tree_mul_77_11_groupi_n_327 & csa_tree_mul_77_11_groupi_n_334)
    | ((csa_tree_mul_77_11_groupi_n_334 & csa_tree_mul_77_11_groupi_n_260) | (csa_tree_mul_77_11_groupi_n_260
    & csa_tree_mul_77_11_groupi_n_327)));
 assign csa_tree_mul_77_11_groupi_n_408 = (csa_tree_mul_77_11_groupi_n_334 ^ (csa_tree_mul_77_11_groupi_n_260
    ^ csa_tree_mul_77_11_groupi_n_327));
 assign csa_tree_mul_77_11_groupi_n_403 = ((csa_tree_mul_77_11_groupi_n_359 & csa_tree_mul_77_11_groupi_n_204)
    | ((csa_tree_mul_77_11_groupi_n_204 & csa_tree_mul_77_11_groupi_n_183) | (csa_tree_mul_77_11_groupi_n_183
    & csa_tree_mul_77_11_groupi_n_359)));
 assign csa_tree_mul_77_11_groupi_n_404 = (csa_tree_mul_77_11_groupi_n_204 ^ (csa_tree_mul_77_11_groupi_n_183
    ^ csa_tree_mul_77_11_groupi_n_359));
 assign csa_tree_mul_77_11_groupi_n_401 = ((csa_tree_mul_77_11_groupi_n_354 & csa_tree_mul_77_11_groupi_n_284)
    | ((csa_tree_mul_77_11_groupi_n_284 & csa_tree_mul_77_11_groupi_n_305) | (csa_tree_mul_77_11_groupi_n_305
    & csa_tree_mul_77_11_groupi_n_354)));
 assign csa_tree_mul_77_11_groupi_n_402 = (csa_tree_mul_77_11_groupi_n_284 ^ (csa_tree_mul_77_11_groupi_n_305
    ^ csa_tree_mul_77_11_groupi_n_354));
 assign csa_tree_mul_77_11_groupi_n_397 = ((csa_tree_mul_77_11_groupi_n_360 & csa_tree_mul_77_11_groupi_n_320)
    | ((csa_tree_mul_77_11_groupi_n_320 & csa_tree_mul_77_11_groupi_n_185) | (csa_tree_mul_77_11_groupi_n_185
    & csa_tree_mul_77_11_groupi_n_360)));
 assign csa_tree_mul_77_11_groupi_n_398 = (csa_tree_mul_77_11_groupi_n_320 ^ (csa_tree_mul_77_11_groupi_n_185
    ^ csa_tree_mul_77_11_groupi_n_360));
 assign csa_tree_mul_77_11_groupi_n_395 = ((csa_tree_mul_77_11_groupi_n_349 & csa_tree_mul_77_11_groupi_n_290)
    | ((csa_tree_mul_77_11_groupi_n_290 & csa_tree_mul_77_11_groupi_n_313) | (csa_tree_mul_77_11_groupi_n_313
    & csa_tree_mul_77_11_groupi_n_349)));
 assign csa_tree_mul_77_11_groupi_n_396 = (csa_tree_mul_77_11_groupi_n_290 ^ (csa_tree_mul_77_11_groupi_n_313
    ^ csa_tree_mul_77_11_groupi_n_349));
 assign csa_tree_mul_77_11_groupi_n_406 = ((csa_tree_mul_77_11_groupi_n_347 & csa_tree_mul_77_11_groupi_n_292)
    | ((csa_tree_mul_77_11_groupi_n_292 & csa_tree_mul_77_11_groupi_n_301) | (csa_tree_mul_77_11_groupi_n_301
    & csa_tree_mul_77_11_groupi_n_347)));
 assign n_1347 = (csa_tree_mul_77_11_groupi_n_292 ^ (csa_tree_mul_77_11_groupi_n_301 ^ csa_tree_mul_77_11_groupi_n_347));
 assign csa_tree_mul_77_11_groupi_n_388 = ((csa_tree_mul_77_11_groupi_n_362 & csa_tree_mul_77_11_groupi_n_282)
    | ((csa_tree_mul_77_11_groupi_n_282 & csa_tree_mul_77_11_groupi_n_182) | (csa_tree_mul_77_11_groupi_n_182
    & csa_tree_mul_77_11_groupi_n_362)));
 assign csa_tree_mul_77_11_groupi_n_389 = (csa_tree_mul_77_11_groupi_n_282 ^ (csa_tree_mul_77_11_groupi_n_182
    ^ csa_tree_mul_77_11_groupi_n_362));
 assign csa_tree_mul_77_11_groupi_n_405 = ~(csa_tree_mul_77_11_groupi_n_384 & csa_tree_mul_77_11_groupi_n_332);
 assign csa_tree_mul_77_11_groupi_n_387 = ~(csa_tree_mul_77_11_groupi_n_384 | csa_tree_mul_77_11_groupi_n_332);
 assign csa_tree_mul_77_11_groupi_n_380 = ((csa_tree_mul_77_11_groupi_n_342 & csa_tree_mul_77_11_groupi_n_280)
    | ((csa_tree_mul_77_11_groupi_n_280 & csa_tree_mul_77_11_groupi_n_210) | (csa_tree_mul_77_11_groupi_n_210
    & csa_tree_mul_77_11_groupi_n_342)));
 assign csa_tree_mul_77_11_groupi_n_381 = (csa_tree_mul_77_11_groupi_n_280 ^ (csa_tree_mul_77_11_groupi_n_210
    ^ csa_tree_mul_77_11_groupi_n_342));
 assign csa_tree_mul_77_11_groupi_n_378 = ((csa_tree_mul_77_11_groupi_n_306 & csa_tree_mul_77_11_groupi_n_309)
    | ((csa_tree_mul_77_11_groupi_n_309 & csa_tree_mul_77_11_groupi_n_203) | (csa_tree_mul_77_11_groupi_n_203
    & csa_tree_mul_77_11_groupi_n_306)));
 assign csa_tree_mul_77_11_groupi_n_379 = (csa_tree_mul_77_11_groupi_n_309 ^ (csa_tree_mul_77_11_groupi_n_203
    ^ csa_tree_mul_77_11_groupi_n_306));
 assign csa_tree_mul_77_11_groupi_n_377 = ((csa_tree_mul_77_11_groupi_n_317 & csa_tree_mul_77_11_groupi_n_201)
    | ((csa_tree_mul_77_11_groupi_n_201 & csa_tree_mul_77_11_groupi_n_197) | (csa_tree_mul_77_11_groupi_n_197
    & csa_tree_mul_77_11_groupi_n_317)));
 assign csa_tree_mul_77_11_groupi_n_385 = (csa_tree_mul_77_11_groupi_n_201 ^ (csa_tree_mul_77_11_groupi_n_197
    ^ csa_tree_mul_77_11_groupi_n_317));
 assign csa_tree_mul_77_11_groupi_n_383 = ((csa_tree_mul_77_11_groupi_n_319 & csa_tree_mul_77_11_groupi_n_289)
    | ((csa_tree_mul_77_11_groupi_n_289 & csa_tree_mul_77_11_groupi_n_195) | (csa_tree_mul_77_11_groupi_n_195
    & csa_tree_mul_77_11_groupi_n_319)));
 assign csa_tree_mul_77_11_groupi_n_384 = (csa_tree_mul_77_11_groupi_n_289 ^ (csa_tree_mul_77_11_groupi_n_195
    ^ csa_tree_mul_77_11_groupi_n_319));
 assign csa_tree_mul_77_11_groupi_n_373 = ((csa_tree_mul_77_11_groupi_n_308 & csa_tree_mul_77_11_groupi_n_202)
    | ((csa_tree_mul_77_11_groupi_n_202 & csa_tree_mul_77_11_groupi_n_184) | (csa_tree_mul_77_11_groupi_n_184
    & csa_tree_mul_77_11_groupi_n_308)));
 assign csa_tree_mul_77_11_groupi_n_374 = (csa_tree_mul_77_11_groupi_n_202 ^ (csa_tree_mul_77_11_groupi_n_184
    ^ csa_tree_mul_77_11_groupi_n_308));
 assign csa_tree_mul_77_11_groupi_n_371 = ((csa_tree_mul_77_11_groupi_n_322 & csa_tree_mul_77_11_groupi_n_283)
    | ((csa_tree_mul_77_11_groupi_n_283 & csa_tree_mul_77_11_groupi_n_199) | (csa_tree_mul_77_11_groupi_n_199
    & csa_tree_mul_77_11_groupi_n_322)));
 assign csa_tree_mul_77_11_groupi_n_372 = (csa_tree_mul_77_11_groupi_n_283 ^ (csa_tree_mul_77_11_groupi_n_199
    ^ csa_tree_mul_77_11_groupi_n_322));
 assign csa_tree_mul_77_11_groupi_n_368 = ((csa_tree_mul_77_11_groupi_n_326 & csa_tree_mul_77_11_groupi_n_287)
    | ((csa_tree_mul_77_11_groupi_n_287 & csa_tree_mul_77_11_groupi_n_247) | (csa_tree_mul_77_11_groupi_n_247
    & csa_tree_mul_77_11_groupi_n_326)));
 assign csa_tree_mul_77_11_groupi_n_369 = (csa_tree_mul_77_11_groupi_n_287 ^ (csa_tree_mul_77_11_groupi_n_247
    ^ csa_tree_mul_77_11_groupi_n_326));
 assign csa_tree_mul_77_11_groupi_n_367 = ~(csa_tree_mul_77_11_groupi_n_344 & csa_tree_mul_77_11_groupi_n_364);
 assign csa_tree_mul_77_11_groupi_n_362 = ((csa_tree_mul_77_11_groupi_n_213 & csa_tree_mul_77_11_groupi_n_223)
    | ((csa_tree_mul_77_11_groupi_n_223 & csa_tree_mul_77_11_groupi_n_259) | (csa_tree_mul_77_11_groupi_n_259
    & csa_tree_mul_77_11_groupi_n_213)));
 assign csa_tree_mul_77_11_groupi_n_363 = (csa_tree_mul_77_11_groupi_n_223 ^ (csa_tree_mul_77_11_groupi_n_259
    ^ csa_tree_mul_77_11_groupi_n_213));
 assign csa_tree_mul_77_11_groupi_n_360 = ((csa_tree_mul_77_11_groupi_n_321 & csa_tree_mul_77_11_groupi_n_288)
    | ((csa_tree_mul_77_11_groupi_n_288 & csa_tree_mul_77_11_groupi_n_189) | (csa_tree_mul_77_11_groupi_n_189
    & csa_tree_mul_77_11_groupi_n_321)));
 assign csa_tree_mul_77_11_groupi_n_361 = (csa_tree_mul_77_11_groupi_n_288 ^ (csa_tree_mul_77_11_groupi_n_189
    ^ csa_tree_mul_77_11_groupi_n_321));
 assign csa_tree_mul_77_11_groupi_n_358 = ((csa_tree_mul_77_11_groupi_n_316 & csa_tree_mul_77_11_groupi_n_257)
    | ((csa_tree_mul_77_11_groupi_n_257 & csa_tree_mul_77_11_groupi_n_158) | (csa_tree_mul_77_11_groupi_n_158
    & csa_tree_mul_77_11_groupi_n_316)));
 assign csa_tree_mul_77_11_groupi_n_359 = (csa_tree_mul_77_11_groupi_n_257 ^ (csa_tree_mul_77_11_groupi_n_158
    ^ csa_tree_mul_77_11_groupi_n_316));
 assign csa_tree_mul_77_11_groupi_n_356 = ((csa_tree_mul_77_11_groupi_n_312 & csa_tree_mul_77_11_groupi_n_196)
    | ((csa_tree_mul_77_11_groupi_n_196 & csa_tree_mul_77_11_groupi_n_200) | (csa_tree_mul_77_11_groupi_n_200
    & csa_tree_mul_77_11_groupi_n_312)));
 assign csa_tree_mul_77_11_groupi_n_357 = (csa_tree_mul_77_11_groupi_n_196 ^ (csa_tree_mul_77_11_groupi_n_200
    ^ csa_tree_mul_77_11_groupi_n_312));
 assign csa_tree_mul_77_11_groupi_n_354 = ((csa_tree_mul_77_11_groupi_n_302 & csa_tree_mul_77_11_groupi_n_190)
    | ((csa_tree_mul_77_11_groupi_n_190 & csa_tree_mul_77_11_groupi_n_193) | (csa_tree_mul_77_11_groupi_n_193
    & csa_tree_mul_77_11_groupi_n_302)));
 assign csa_tree_mul_77_11_groupi_n_355 = (csa_tree_mul_77_11_groupi_n_190 ^ (csa_tree_mul_77_11_groupi_n_193
    ^ csa_tree_mul_77_11_groupi_n_302));
 assign csa_tree_mul_77_11_groupi_n_352 = (csa_tree_mul_77_11_groupi_n_307 & csa_tree_mul_77_11_groupi_n_214);
 assign csa_tree_mul_77_11_groupi_n_353 = (csa_tree_mul_77_11_groupi_n_307 ^ csa_tree_mul_77_11_groupi_n_214);
 assign csa_tree_mul_77_11_groupi_n_365 = ((csa_tree_mul_77_11_groupi_n_318 & csa_tree_mul_77_11_groupi_n_198)
    | ((csa_tree_mul_77_11_groupi_n_198 & csa_tree_mul_77_11_groupi_n_173) | (csa_tree_mul_77_11_groupi_n_173
    & csa_tree_mul_77_11_groupi_n_318)));
 assign csa_tree_mul_77_11_groupi_n_351 = (csa_tree_mul_77_11_groupi_n_198 ^ (csa_tree_mul_77_11_groupi_n_173
    ^ csa_tree_mul_77_11_groupi_n_318));
 assign csa_tree_mul_77_11_groupi_n_349 = ((csa_tree_mul_77_11_groupi_n_303 & csa_tree_mul_77_11_groupi_n_278)
    | ((csa_tree_mul_77_11_groupi_n_278 & csa_tree_mul_77_11_groupi_n_207) | (csa_tree_mul_77_11_groupi_n_207
    & csa_tree_mul_77_11_groupi_n_303)));
 assign csa_tree_mul_77_11_groupi_n_350 = (csa_tree_mul_77_11_groupi_n_278 ^ (csa_tree_mul_77_11_groupi_n_207
    ^ csa_tree_mul_77_11_groupi_n_303));
 assign csa_tree_mul_77_11_groupi_n_347 = ((csa_tree_mul_77_11_groupi_n_314 & csa_tree_mul_77_11_groupi_n_294)
    | ((csa_tree_mul_77_11_groupi_n_294 & csa_tree_mul_77_11_groupi_n_160) | (csa_tree_mul_77_11_groupi_n_160
    & csa_tree_mul_77_11_groupi_n_314)));
 assign n_1348 = (csa_tree_mul_77_11_groupi_n_294 ^ (csa_tree_mul_77_11_groupi_n_160 ^ csa_tree_mul_77_11_groupi_n_314));
 assign csa_tree_mul_77_11_groupi_n_345 = ((csa_tree_mul_77_11_groupi_n_325 & csa_tree_mul_77_11_groupi_n_187)
    | ((csa_tree_mul_77_11_groupi_n_187 & csa_tree_mul_77_11_groupi_n_194) | (csa_tree_mul_77_11_groupi_n_194
    & csa_tree_mul_77_11_groupi_n_325)));
 assign csa_tree_mul_77_11_groupi_n_346 = (csa_tree_mul_77_11_groupi_n_187 ^ (csa_tree_mul_77_11_groupi_n_194
    ^ csa_tree_mul_77_11_groupi_n_325));
 assign csa_tree_mul_77_11_groupi_n_364 = ~(csa_tree_mul_77_11_groupi_n_333 & csa_tree_mul_77_11_groupi_n_296);
 assign csa_tree_mul_77_11_groupi_n_344 = (csa_tree_mul_77_11_groupi_n_333 | csa_tree_mul_77_11_groupi_n_296);
 assign csa_tree_mul_77_11_groupi_n_342 = ((csa_tree_mul_77_11_groupi_n_232 & csa_tree_mul_77_11_groupi_n_188)
    | ((csa_tree_mul_77_11_groupi_n_188 & csa_tree_mul_77_11_groupi_n_262) | (csa_tree_mul_77_11_groupi_n_262
    & csa_tree_mul_77_11_groupi_n_232)));
 assign csa_tree_mul_77_11_groupi_n_343 = (csa_tree_mul_77_11_groupi_n_188 ^ (csa_tree_mul_77_11_groupi_n_262
    ^ csa_tree_mul_77_11_groupi_n_232));
 assign csa_tree_mul_77_11_groupi_n_338 = ((csa_tree_mul_77_11_groupi_n_227 & csa_tree_mul_77_11_groupi_n_186)
    | ((csa_tree_mul_77_11_groupi_n_186 & csa_tree_mul_77_11_groupi_n_258) | (csa_tree_mul_77_11_groupi_n_258
    & csa_tree_mul_77_11_groupi_n_227)));
 assign csa_tree_mul_77_11_groupi_n_339 = (csa_tree_mul_77_11_groupi_n_186 ^ (csa_tree_mul_77_11_groupi_n_258
    ^ csa_tree_mul_77_11_groupi_n_227));
 assign csa_tree_mul_77_11_groupi_n_334 = ((csa_tree_mul_77_11_groupi_n_251 & csa_tree_mul_77_11_groupi_n_218)
    | ((csa_tree_mul_77_11_groupi_n_218 & csa_tree_mul_77_11_groupi_n_261) | (csa_tree_mul_77_11_groupi_n_261
    & csa_tree_mul_77_11_groupi_n_251)));
 assign csa_tree_mul_77_11_groupi_n_335 = (csa_tree_mul_77_11_groupi_n_218 ^ (csa_tree_mul_77_11_groupi_n_261
    ^ csa_tree_mul_77_11_groupi_n_251));
 assign csa_tree_mul_77_11_groupi_n_332 = ((csa_tree_mul_77_11_groupi_n_300 & csa_tree_mul_77_11_groupi_n_222)
    | ((csa_tree_mul_77_11_groupi_n_222 & csa_tree_mul_77_11_groupi_n_159) | (csa_tree_mul_77_11_groupi_n_159
    & csa_tree_mul_77_11_groupi_n_300)));
 assign csa_tree_mul_77_11_groupi_n_333 = (csa_tree_mul_77_11_groupi_n_222 ^ (csa_tree_mul_77_11_groupi_n_159
    ^ csa_tree_mul_77_11_groupi_n_300));
 assign csa_tree_mul_77_11_groupi_n_330 = ((csa_tree_mul_77_11_groupi_n_273 & csa_tree_mul_77_11_groupi_n_219)
    | ((csa_tree_mul_77_11_groupi_n_219 & csa_tree_mul_77_11_groupi_n_226) | (csa_tree_mul_77_11_groupi_n_226
    & csa_tree_mul_77_11_groupi_n_273)));
 assign csa_tree_mul_77_11_groupi_n_331 = (csa_tree_mul_77_11_groupi_n_219 ^ (csa_tree_mul_77_11_groupi_n_226
    ^ csa_tree_mul_77_11_groupi_n_273));
 assign csa_tree_mul_77_11_groupi_n_328 = ((csa_tree_mul_77_11_groupi_n_291 & csa_tree_mul_77_11_groupi_n_221)
    | ((csa_tree_mul_77_11_groupi_n_221 & csa_tree_mul_77_11_groupi_n_248) | (csa_tree_mul_77_11_groupi_n_248
    & csa_tree_mul_77_11_groupi_n_291)));
 assign csa_tree_mul_77_11_groupi_n_329 = (csa_tree_mul_77_11_groupi_n_221 ^ (csa_tree_mul_77_11_groupi_n_248
    ^ csa_tree_mul_77_11_groupi_n_291));
 assign csa_tree_mul_77_11_groupi_n_326 = ((csa_tree_mul_77_11_groupi_n_237 & csa_tree_mul_77_11_groupi_n_252)
    | ((csa_tree_mul_77_11_groupi_n_252 & csa_tree_mul_77_11_groupi_n_217) | (csa_tree_mul_77_11_groupi_n_217
    & csa_tree_mul_77_11_groupi_n_237)));
 assign csa_tree_mul_77_11_groupi_n_327 = (csa_tree_mul_77_11_groupi_n_252 ^ (csa_tree_mul_77_11_groupi_n_217
    ^ csa_tree_mul_77_11_groupi_n_237));
 assign csa_tree_mul_77_11_groupi_n_324 = (csa_tree_mul_77_11_groupi_n_271 & csa_tree_mul_77_11_groupi_n_229);
 assign csa_tree_mul_77_11_groupi_n_325 = (csa_tree_mul_77_11_groupi_n_271 ^ csa_tree_mul_77_11_groupi_n_229);
 assign csa_tree_mul_77_11_groupi_n_322 = (csa_tree_mul_77_11_groupi_n_268 & csa_tree_mul_77_11_groupi_n_233);
 assign csa_tree_mul_77_11_groupi_n_323 = (csa_tree_mul_77_11_groupi_n_268 ^ csa_tree_mul_77_11_groupi_n_233);
 assign csa_tree_mul_77_11_groupi_n_320 = (csa_tree_mul_77_11_groupi_n_267 & csa_tree_mul_77_11_groupi_n_236);
 assign csa_tree_mul_77_11_groupi_n_321 = (csa_tree_mul_77_11_groupi_n_267 ^ csa_tree_mul_77_11_groupi_n_236);
 assign csa_tree_mul_77_11_groupi_n_318 = (csa_tree_mul_77_11_groupi_n_216 & csa_tree_mul_77_11_groupi_n_263);
 assign csa_tree_mul_77_11_groupi_n_319 = (csa_tree_mul_77_11_groupi_n_216 ^ csa_tree_mul_77_11_groupi_n_263);
 assign csa_tree_mul_77_11_groupi_n_316 = (csa_tree_mul_77_11_groupi_n_265 & csa_tree_mul_77_11_groupi_n_275);
 assign csa_tree_mul_77_11_groupi_n_317 = (csa_tree_mul_77_11_groupi_n_265 ^ csa_tree_mul_77_11_groupi_n_275);
 assign csa_tree_mul_77_11_groupi_n_314 = (csa_tree_mul_77_11_groupi_n_293 & csa_tree_mul_77_11_groupi_n_98);
 assign n_1349 = (csa_tree_mul_77_11_groupi_n_293 ^ csa_tree_mul_77_11_groupi_n_98);
 assign csa_tree_mul_77_11_groupi_n_312 = (csa_tree_mul_77_11_groupi_n_272 & csa_tree_mul_77_11_groupi_n_238);
 assign csa_tree_mul_77_11_groupi_n_313 = (csa_tree_mul_77_11_groupi_n_272 ^ csa_tree_mul_77_11_groupi_n_238);
 assign csa_tree_mul_77_11_groupi_n_310 = (csa_tree_mul_77_11_groupi_n_269 & csa_tree_mul_77_11_groupi_n_234);
 assign csa_tree_mul_77_11_groupi_n_311 = (csa_tree_mul_77_11_groupi_n_269 ^ csa_tree_mul_77_11_groupi_n_234);
 assign csa_tree_mul_77_11_groupi_n_308 = (csa_tree_mul_77_11_groupi_n_274 & csa_tree_mul_77_11_groupi_n_235);
 assign csa_tree_mul_77_11_groupi_n_309 = (csa_tree_mul_77_11_groupi_n_274 ^ csa_tree_mul_77_11_groupi_n_235);
 assign csa_tree_mul_77_11_groupi_n_306 = (csa_tree_mul_77_11_groupi_n_264 & csa_tree_mul_77_11_groupi_n_228);
 assign csa_tree_mul_77_11_groupi_n_307 = (csa_tree_mul_77_11_groupi_n_264 ^ csa_tree_mul_77_11_groupi_n_228);
 assign csa_tree_mul_77_11_groupi_n_304 = (csa_tree_mul_77_11_groupi_n_270 & csa_tree_mul_77_11_groupi_n_230);
 assign csa_tree_mul_77_11_groupi_n_305 = (csa_tree_mul_77_11_groupi_n_270 ^ csa_tree_mul_77_11_groupi_n_230);
 assign csa_tree_mul_77_11_groupi_n_302 = (csa_tree_mul_77_11_groupi_n_266 & csa_tree_mul_77_11_groupi_n_231);
 assign csa_tree_mul_77_11_groupi_n_303 = (csa_tree_mul_77_11_groupi_n_266 ^ csa_tree_mul_77_11_groupi_n_231);
 assign csa_tree_mul_77_11_groupi_n_300 = (csa_tree_mul_77_11_groupi_n_211 & csa_tree_mul_77_11_groupi_n_166);
 assign csa_tree_mul_77_11_groupi_n_301 = (csa_tree_mul_77_11_groupi_n_211 ^ csa_tree_mul_77_11_groupi_n_166);
 assign csa_tree_mul_77_11_groupi_n_299 = ~(csa_tree_mul_77_11_groupi_n_298 & (csa_tree_mul_77_11_groupi_n_253
    | csa_tree_mul_77_11_groupi_n_297));
 assign csa_tree_mul_77_11_groupi_n_298 = ~(csa_tree_mul_77_11_groupi_n_253 & csa_tree_mul_77_11_groupi_n_297);
 assign csa_tree_mul_77_11_groupi_n_297 = ~(csa_tree_mul_77_11_groupi_n_39 & ~(csa_tree_mul_77_11_groupi_n_178
    & n_1321));
 assign csa_tree_mul_77_11_groupi_n_294 = ~((n_1489 | csa_tree_mul_77_11_groupi_n_96) & (csa_tree_mul_77_11_groupi_n_85
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_296 = ~((n_1489 | csa_tree_mul_77_11_groupi_n_81) & (csa_tree_mul_77_11_groupi_n_95
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_293 = ~((n_1489 | csa_tree_mul_77_11_groupi_n_52) & (csa_tree_mul_77_11_groupi_n_96
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_292 = ~((n_1489 | csa_tree_mul_77_11_groupi_n_85) & (csa_tree_mul_77_11_groupi_n_81
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_291 = ~(csa_tree_mul_77_11_groupi_n_181 | (csa_tree_mul_77_11_groupi_n_176
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_290 = ~((n_1489 | csa_tree_mul_77_11_groupi_n_86) & (csa_tree_mul_77_11_groupi_n_91
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_289 = ~(csa_tree_mul_77_11_groupi_n_244 & (csa_tree_mul_77_11_groupi_n_84
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_288 = ~((n_1489 | csa_tree_mul_77_11_groupi_n_93) & (csa_tree_mul_77_11_groupi_n_94
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_287 = ~(csa_tree_mul_77_11_groupi_n_180 & ~(csa_tree_mul_77_11_groupi_n_176
    & csa_tree_mul_77_11_groupi_n_64));
 assign csa_tree_mul_77_11_groupi_n_286 = ~(csa_tree_mul_77_11_groupi_n_245 & (csa_tree_mul_77_11_groupi_n_88
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_285 = ~(csa_tree_mul_77_11_groupi_n_39 & ~(csa_tree_mul_77_11_groupi_n_178
    & csa_tree_mul_77_11_groupi_n_90));
 assign csa_tree_mul_77_11_groupi_n_284 = ~((n_1489 | csa_tree_mul_77_11_groupi_n_91) & (csa_tree_mul_77_11_groupi_n_89
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_295 = ~(csa_tree_mul_77_11_groupi_n_1 & (n_1491 | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_283 = ~(csa_tree_mul_77_11_groupi_n_246 & (csa_tree_mul_77_11_groupi_n_93
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_282 = ~((n_1489 | csa_tree_mul_77_11_groupi_n_55) & (csa_tree_mul_77_11_groupi_n_87
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_281 = ~(csa_tree_mul_77_11_groupi_n_239 & (csa_tree_mul_77_11_groupi_n_92
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_280 = ~((n_1489 | csa_tree_mul_77_11_groupi_n_83) & (csa_tree_mul_77_11_groupi_n_55
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_279 = ~(csa_tree_mul_77_11_groupi_n_243 & ~(csa_tree_mul_77_11_groupi_n_82
    & n_1322));
 assign csa_tree_mul_77_11_groupi_n_278 = ~((n_1489 | csa_tree_mul_77_11_groupi_n_94) & (csa_tree_mul_77_11_groupi_n_86
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_277 = ~(csa_tree_mul_77_11_groupi_n_241 & (csa_tree_mul_77_11_groupi_n_97
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_276 = ~((n_1489 | csa_tree_mul_77_11_groupi_n_88) & (csa_tree_mul_77_11_groupi_n_54
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_275 = ~(csa_tree_mul_77_11_groupi_n_28 | ((csa_tree_mul_77_11_groupi_n_47
    & n_1313) | (n_1317 & n_1316)));
 assign csa_tree_mul_77_11_groupi_n_274 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_62)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_78));
 assign csa_tree_mul_77_11_groupi_n_273 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_79)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_77));
 assign csa_tree_mul_77_11_groupi_n_272 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_68)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_65));
 assign csa_tree_mul_77_11_groupi_n_271 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_72)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_70));
 assign csa_tree_mul_77_11_groupi_n_270 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_65)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_72));
 assign csa_tree_mul_77_11_groupi_n_269 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_69)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_67));
 assign csa_tree_mul_77_11_groupi_n_268 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_78)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_69));
 assign csa_tree_mul_77_11_groupi_n_267 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_67)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_76));
 assign csa_tree_mul_77_11_groupi_n_266 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_76)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_68));
 assign csa_tree_mul_77_11_groupi_n_265 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_49)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_66));
 assign csa_tree_mul_77_11_groupi_n_264 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_61)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_62));
 assign csa_tree_mul_77_11_groupi_n_263 = ~(csa_tree_mul_77_11_groupi_n_27 | ((n_1319 & n_1313) | (csa_tree_mul_77_11_groupi_n_40
    & n_1318)));
 assign csa_tree_mul_77_11_groupi_n_262 = ~(csa_tree_mul_77_11_groupi_n_240 & ~(csa_tree_mul_77_11_groupi_n_165
    & csa_tree_mul_77_11_groupi_n_74));
 assign csa_tree_mul_77_11_groupi_n_261 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_77)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_59));
 assign csa_tree_mul_77_11_groupi_n_260 = ((csa_tree_mul_77_11_groupi_n_165 & csa_tree_mul_77_11_groupi_n_64)
    | (csa_tree_mul_77_11_groupi_n_176 & csa_tree_mul_77_11_groupi_n_60));
 assign csa_tree_mul_77_11_groupi_n_259 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_75)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_61));
 assign csa_tree_mul_77_11_groupi_n_258 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_73)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_71));
 assign csa_tree_mul_77_11_groupi_n_257 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_66)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_73));
 assign csa_tree_mul_77_11_groupi_n_256 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_63)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_79));
 assign csa_tree_mul_77_11_groupi_n_255 = ~(csa_tree_mul_77_11_groupi_n_242 & (csa_tree_mul_77_11_groupi_n_80
    | csa_tree_mul_77_11_groupi_n_14));
 assign csa_tree_mul_77_11_groupi_n_254 = ~((csa_tree_mul_77_11_groupi_n_177 | csa_tree_mul_77_11_groupi_n_70)
    & (csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_63));
 assign csa_tree_mul_77_11_groupi_n_252 = ~csa_tree_mul_77_11_groupi_n_251;
 assign csa_tree_mul_77_11_groupi_n_250 = ~csa_tree_mul_77_11_groupi_n_249;
 assign csa_tree_mul_77_11_groupi_n_248 = ~csa_tree_mul_77_11_groupi_n_247;
 assign csa_tree_mul_77_11_groupi_n_246 = ~(csa_tree_mul_77_11_groupi_n_178 & ~csa_tree_mul_77_11_groupi_n_54);
 assign csa_tree_mul_77_11_groupi_n_245 = ~(csa_tree_mul_77_11_groupi_n_178 & ~csa_tree_mul_77_11_groupi_n_87);
 assign csa_tree_mul_77_11_groupi_n_244 = ~(csa_tree_mul_77_11_groupi_n_178 & ~csa_tree_mul_77_11_groupi_n_95);
 assign csa_tree_mul_77_11_groupi_n_243 = ~(csa_tree_mul_77_11_groupi_n_178 & ~csa_tree_mul_77_11_groupi_n_97);
 assign csa_tree_mul_77_11_groupi_n_242 = ~(csa_tree_mul_77_11_groupi_n_178 & ~n_1491);
 assign csa_tree_mul_77_11_groupi_n_241 = ~(csa_tree_mul_77_11_groupi_n_178 & ~csa_tree_mul_77_11_groupi_n_80);
 assign csa_tree_mul_77_11_groupi_n_240 = ~(csa_tree_mul_77_11_groupi_n_176 & ~csa_tree_mul_77_11_groupi_n_71);
 assign csa_tree_mul_77_11_groupi_n_239 = ~(csa_tree_mul_77_11_groupi_n_178 & ~csa_tree_mul_77_11_groupi_n_84);
 assign csa_tree_mul_77_11_groupi_n_253 = ~((csa_tree_mul_77_11_groupi_n_163 & n_1301) | (csa_tree_mul_77_11_groupi_n_107
    & n_1300));
 assign csa_tree_mul_77_11_groupi_n_238 = ~((csa_tree_mul_77_11_groupi_n_164 | csa_tree_mul_77_11_groupi_n_25)
    & (csa_tree_mul_77_11_groupi_n_0 | csa_tree_mul_77_11_groupi_n_36));
 assign csa_tree_mul_77_11_groupi_n_237 = ~((csa_tree_mul_77_11_groupi_n_164 | csa_tree_mul_77_11_groupi_n_35)
    & (csa_tree_mul_77_11_groupi_n_0 | csa_tree_mul_77_11_groupi_n_31));
 assign csa_tree_mul_77_11_groupi_n_236 = ~((csa_tree_mul_77_11_groupi_n_164 | csa_tree_mul_77_11_groupi_n_16)
    & (csa_tree_mul_77_11_groupi_n_0 | csa_tree_mul_77_11_groupi_n_21));
 assign csa_tree_mul_77_11_groupi_n_235 = ~((csa_tree_mul_77_11_groupi_n_164 | csa_tree_mul_77_11_groupi_n_19)
    & (csa_tree_mul_77_11_groupi_n_0 | csa_tree_mul_77_11_groupi_n_20));
 assign csa_tree_mul_77_11_groupi_n_234 = ~((csa_tree_mul_77_11_groupi_n_164 | csa_tree_mul_77_11_groupi_n_33)
    & (csa_tree_mul_77_11_groupi_n_0 | csa_tree_mul_77_11_groupi_n_16));
 assign csa_tree_mul_77_11_groupi_n_233 = ~((csa_tree_mul_77_11_groupi_n_164 | csa_tree_mul_77_11_groupi_n_20)
    & (csa_tree_mul_77_11_groupi_n_0 | csa_tree_mul_77_11_groupi_n_33));
 assign csa_tree_mul_77_11_groupi_n_232 = ~((csa_tree_mul_77_11_groupi_n_164 | csa_tree_mul_77_11_groupi_n_22)
    & (csa_tree_mul_77_11_groupi_n_0 | csa_tree_mul_77_11_groupi_n_37));
 assign csa_tree_mul_77_11_groupi_n_231 = ~((csa_tree_mul_77_11_groupi_n_164 | csa_tree_mul_77_11_groupi_n_21)
    & (csa_tree_mul_77_11_groupi_n_0 | csa_tree_mul_77_11_groupi_n_25));
 assign csa_tree_mul_77_11_groupi_n_230 = ~((csa_tree_mul_77_11_groupi_n_164 | csa_tree_mul_77_11_groupi_n_36)
    & (csa_tree_mul_77_11_groupi_n_0 | csa_tree_mul_77_11_groupi_n_18));
 assign csa_tree_mul_77_11_groupi_n_229 = ~((csa_tree_mul_77_11_groupi_n_164 | csa_tree_mul_77_11_groupi_n_18)
    & (csa_tree_mul_77_11_groupi_n_0 | csa_tree_mul_77_11_groupi_n_34));
 assign csa_tree_mul_77_11_groupi_n_228 = ~((csa_tree_mul_77_11_groupi_n_164 | csa_tree_mul_77_11_groupi_n_23)
    & (csa_tree_mul_77_11_groupi_n_0 | csa_tree_mul_77_11_groupi_n_19));
 assign csa_tree_mul_77_11_groupi_n_227 = ~((csa_tree_mul_77_11_groupi_n_164 | csa_tree_mul_77_11_groupi_n_29)
    & (csa_tree_mul_77_11_groupi_n_0 | csa_tree_mul_77_11_groupi_n_22));
 assign csa_tree_mul_77_11_groupi_n_226 = ~(csa_tree_mul_77_11_groupi_n_155 | (csa_tree_mul_77_11_groupi_n_162
    & n_1319));
 assign csa_tree_mul_77_11_groupi_n_225 = ~((csa_tree_mul_77_11_groupi_n_161 | csa_tree_mul_77_11_groupi_n_126)
    & (csa_tree_mul_77_11_groupi_n_106 | csa_tree_mul_77_11_groupi_n_121));
 assign csa_tree_mul_77_11_groupi_n_224 = ~(csa_tree_mul_77_11_groupi_n_154 & ~(csa_tree_mul_77_11_groupi_n_162
    & csa_tree_mul_77_11_groupi_n_122));
 assign csa_tree_mul_77_11_groupi_n_223 = ~((csa_tree_mul_77_11_groupi_n_164 | csa_tree_mul_77_11_groupi_n_37)
    & (csa_tree_mul_77_11_groupi_n_0 | csa_tree_mul_77_11_groupi_n_23));
 assign csa_tree_mul_77_11_groupi_n_222 = ~((csa_tree_mul_77_11_groupi_n_161 | csa_tree_mul_77_11_groupi_n_133)
    & (csa_tree_mul_77_11_groupi_n_106 | csa_tree_mul_77_11_groupi_n_148));
 assign csa_tree_mul_77_11_groupi_n_221 = ~((csa_tree_mul_77_11_groupi_n_164 | csa_tree_mul_77_11_groupi_n_17)
    & (csa_tree_mul_77_11_groupi_n_0 | csa_tree_mul_77_11_groupi_n_30));
 assign csa_tree_mul_77_11_groupi_n_220 = ~(csa_tree_mul_77_11_groupi_n_172 & ~(csa_tree_mul_77_11_groupi_n_105
    & csa_tree_mul_77_11_groupi_n_145));
 assign csa_tree_mul_77_11_groupi_n_219 = ~((csa_tree_mul_77_11_groupi_n_164 | csa_tree_mul_77_11_groupi_n_24)
    & (csa_tree_mul_77_11_groupi_n_0 | csa_tree_mul_77_11_groupi_n_32));
 assign csa_tree_mul_77_11_groupi_n_218 = ~(csa_tree_mul_77_11_groupi_n_156 & ~(csa_tree_mul_77_11_groupi_n_152
    & csa_tree_mul_77_11_groupi_n_117));
 assign csa_tree_mul_77_11_groupi_n_217 = ~(csa_tree_mul_77_11_groupi_n_157 | (csa_tree_mul_77_11_groupi_n_152
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_251 = ~((csa_tree_mul_77_11_groupi_n_163 & n_1298) | (csa_tree_mul_77_11_groupi_n_107
    & n_1297));
 assign csa_tree_mul_77_11_groupi_n_249 = ~((csa_tree_mul_77_11_groupi_n_163 & n_1300) | (csa_tree_mul_77_11_groupi_n_107
    & n_1299));
 assign csa_tree_mul_77_11_groupi_n_247 = ~((csa_tree_mul_77_11_groupi_n_163 & n_1296) | (csa_tree_mul_77_11_groupi_n_107
    & n_1295));
 assign csa_tree_mul_77_11_groupi_n_216 = ~((csa_tree_mul_77_11_groupi_n_153 | csa_tree_mul_77_11_groupi_n_50)
    & (csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_129));
 assign csa_tree_mul_77_11_groupi_n_215 = ~((csa_tree_mul_77_11_groupi_n_153 | csa_tree_mul_77_11_groupi_n_132)
    & (csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_115));
 assign csa_tree_mul_77_11_groupi_n_214 = ~((csa_tree_mul_77_11_groupi_n_153 | csa_tree_mul_77_11_groupi_n_141)
    & (csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_120));
 assign csa_tree_mul_77_11_groupi_n_213 = ~((csa_tree_mul_77_11_groupi_n_153 | csa_tree_mul_77_11_groupi_n_137)
    & (csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_141));
 assign csa_tree_mul_77_11_groupi_n_212 = ~((csa_tree_mul_77_11_groupi_n_153 | csa_tree_mul_77_11_groupi_n_115)
    & (csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_110));
 assign csa_tree_mul_77_11_groupi_n_211 = ~((csa_tree_mul_77_11_groupi_n_161 | csa_tree_mul_77_11_groupi_n_51)
    & (csa_tree_mul_77_11_groupi_n_106 | csa_tree_mul_77_11_groupi_n_133));
 assign csa_tree_mul_77_11_groupi_n_210 = ~(csa_tree_mul_77_11_groupi_n_150 & ~(csa_tree_mul_77_11_groupi_n_162
    & csa_tree_mul_77_11_groupi_n_109));
 assign csa_tree_mul_77_11_groupi_n_209 = ~((csa_tree_mul_77_11_groupi_n_161 | csa_tree_mul_77_11_groupi_n_121)
    & (csa_tree_mul_77_11_groupi_n_106 | csa_tree_mul_77_11_groupi_n_123));
 assign csa_tree_mul_77_11_groupi_n_208 = ~(csa_tree_mul_77_11_groupi_n_170 & (csa_tree_mul_77_11_groupi_n_106
    | n_1490));
 assign csa_tree_mul_77_11_groupi_n_207 = ~((csa_tree_mul_77_11_groupi_n_161 | csa_tree_mul_77_11_groupi_n_123)
    & (csa_tree_mul_77_11_groupi_n_106 | csa_tree_mul_77_11_groupi_n_114));
 assign csa_tree_mul_77_11_groupi_n_206 = ~(csa_tree_mul_77_11_groupi_n_169 & ~(csa_tree_mul_77_11_groupi_n_105
    & csa_tree_mul_77_11_groupi_n_128));
 assign csa_tree_mul_77_11_groupi_n_205 = ((csa_tree_mul_77_11_groupi_n_105 & csa_tree_mul_77_11_groupi_n_122)
    | (csa_tree_mul_77_11_groupi_n_162 & csa_tree_mul_77_11_groupi_n_119));
 assign csa_tree_mul_77_11_groupi_n_204 = ~(csa_tree_mul_77_11_groupi_n_168 & ~(csa_tree_mul_77_11_groupi_n_105
    & csa_tree_mul_77_11_groupi_n_131));
 assign csa_tree_mul_77_11_groupi_n_203 = ~((csa_tree_mul_77_11_groupi_n_161 | csa_tree_mul_77_11_groupi_n_113)
    & (csa_tree_mul_77_11_groupi_n_106 | csa_tree_mul_77_11_groupi_n_142));
 assign csa_tree_mul_77_11_groupi_n_202 = ~(csa_tree_mul_77_11_groupi_n_151 & ~(csa_tree_mul_77_11_groupi_n_162
    & csa_tree_mul_77_11_groupi_n_143));
 assign csa_tree_mul_77_11_groupi_n_201 = ~(csa_tree_mul_77_11_groupi_n_171 & (csa_tree_mul_77_11_groupi_n_106
    | csa_tree_mul_77_11_groupi_n_135));
 assign csa_tree_mul_77_11_groupi_n_200 = ~((csa_tree_mul_77_11_groupi_n_153 | csa_tree_mul_77_11_groupi_n_130)
    & (csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_116));
 assign csa_tree_mul_77_11_groupi_n_199 = ~((csa_tree_mul_77_11_groupi_n_153 | csa_tree_mul_77_11_groupi_n_124)
    & (csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_112));
 assign csa_tree_mul_77_11_groupi_n_198 = ~((csa_tree_mul_77_11_groupi_n_153 | csa_tree_mul_77_11_groupi_n_129)
    & (csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_138));
 assign csa_tree_mul_77_11_groupi_n_197 = ~((csa_tree_mul_77_11_groupi_n_153 | csa_tree_mul_77_11_groupi_n_138)
    & (csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_146));
 assign csa_tree_mul_77_11_groupi_n_196 = ~((csa_tree_mul_77_11_groupi_n_161 | csa_tree_mul_77_11_groupi_n_147)
    & (csa_tree_mul_77_11_groupi_n_106 | csa_tree_mul_77_11_groupi_n_140));
 assign csa_tree_mul_77_11_groupi_n_195 = ~((csa_tree_mul_77_11_groupi_n_161 | csa_tree_mul_77_11_groupi_n_148)
    & (csa_tree_mul_77_11_groupi_n_106 | csa_tree_mul_77_11_groupi_n_127));
 assign csa_tree_mul_77_11_groupi_n_194 = ~((csa_tree_mul_77_11_groupi_n_153 | csa_tree_mul_77_11_groupi_n_116)
    & (csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_132));
 assign csa_tree_mul_77_11_groupi_n_193 = ~((csa_tree_mul_77_11_groupi_n_153 | csa_tree_mul_77_11_groupi_n_58)
    & (csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_130));
 assign csa_tree_mul_77_11_groupi_n_192 = ((csa_tree_mul_77_11_groupi_n_102 & csa_tree_mul_77_11_groupi_n_117)
    | (csa_tree_mul_77_11_groupi_n_152 & csa_tree_mul_77_11_groupi_n_111));
 assign csa_tree_mul_77_11_groupi_n_191 = ~((csa_tree_mul_77_11_groupi_n_153 | csa_tree_mul_77_11_groupi_n_120)
    & (csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_149));
 assign csa_tree_mul_77_11_groupi_n_190 = ~((csa_tree_mul_77_11_groupi_n_161 | csa_tree_mul_77_11_groupi_n_114)
    & (csa_tree_mul_77_11_groupi_n_106 | csa_tree_mul_77_11_groupi_n_147));
 assign csa_tree_mul_77_11_groupi_n_189 = ~((csa_tree_mul_77_11_groupi_n_153 | csa_tree_mul_77_11_groupi_n_112)
    & (csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_139));
 assign csa_tree_mul_77_11_groupi_n_188 = ~(csa_tree_mul_77_11_groupi_n_175 & ~(csa_tree_mul_77_11_groupi_n_102
    & csa_tree_mul_77_11_groupi_n_136));
 assign csa_tree_mul_77_11_groupi_n_187 = ~((csa_tree_mul_77_11_groupi_n_161 | csa_tree_mul_77_11_groupi_n_140)
    & (csa_tree_mul_77_11_groupi_n_106 | csa_tree_mul_77_11_groupi_n_118));
 assign csa_tree_mul_77_11_groupi_n_186 = ~(csa_tree_mul_77_11_groupi_n_167 & (csa_tree_mul_77_11_groupi_n_103
    | csa_tree_mul_77_11_groupi_n_134));
 assign csa_tree_mul_77_11_groupi_n_185 = ~((csa_tree_mul_77_11_groupi_n_153 | csa_tree_mul_77_11_groupi_n_139)
    & (csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_58));
 assign csa_tree_mul_77_11_groupi_n_184 = ~((csa_tree_mul_77_11_groupi_n_153 | csa_tree_mul_77_11_groupi_n_149)
    & (csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_124));
 assign csa_tree_mul_77_11_groupi_n_183 = ~((csa_tree_mul_77_11_groupi_n_153 | csa_tree_mul_77_11_groupi_n_146)
    & (csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_144));
 assign csa_tree_mul_77_11_groupi_n_182 = ~((csa_tree_mul_77_11_groupi_n_161 | csa_tree_mul_77_11_groupi_n_57)
    & (csa_tree_mul_77_11_groupi_n_106 | csa_tree_mul_77_11_groupi_n_113));
 assign csa_tree_mul_77_11_groupi_n_181 = ~csa_tree_mul_77_11_groupi_n_180;
 assign csa_tree_mul_77_11_groupi_n_178 = ~n_1489;
 assign csa_tree_mul_77_11_groupi_n_176 = ~csa_tree_mul_77_11_groupi_n_177;
 assign csa_tree_mul_77_11_groupi_n_175 = ~(csa_tree_mul_77_11_groupi_n_152 & ~csa_tree_mul_77_11_groupi_n_134);
 assign csa_tree_mul_77_11_groupi_n_174 = ~(csa_tree_mul_77_11_groupi_n_164 | csa_tree_mul_77_11_groupi_n_30);
 assign csa_tree_mul_77_11_groupi_n_180 = ~(csa_tree_mul_77_11_groupi_n_165 & n_1315);
 assign csa_tree_mul_77_11_groupi_n_173 = ~(csa_tree_mul_77_11_groupi_n_104 | csa_tree_mul_77_11_groupi_n_29);
 assign csa_tree_mul_77_11_groupi_n_177 = (csa_tree_mul_77_11_groupi_n_165 | csa_tree_mul_77_11_groupi_n_99);
 assign csa_tree_mul_77_11_groupi_n_172 = ~(csa_tree_mul_77_11_groupi_n_162 & ~csa_tree_mul_77_11_groupi_n_127);
 assign csa_tree_mul_77_11_groupi_n_171 = ~(csa_tree_mul_77_11_groupi_n_162 & csa_tree_mul_77_11_groupi_n_145);
 assign csa_tree_mul_77_11_groupi_n_170 = ~(csa_tree_mul_77_11_groupi_n_128 & ~csa_tree_mul_77_11_groupi_n_161);
 assign csa_tree_mul_77_11_groupi_n_169 = ~(csa_tree_mul_77_11_groupi_n_131 & ~csa_tree_mul_77_11_groupi_n_161);
 assign csa_tree_mul_77_11_groupi_n_168 = ~(csa_tree_mul_77_11_groupi_n_162 & ~csa_tree_mul_77_11_groupi_n_135);
 assign csa_tree_mul_77_11_groupi_n_167 = ~(csa_tree_mul_77_11_groupi_n_152 & ~csa_tree_mul_77_11_groupi_n_144);
 assign csa_tree_mul_77_11_groupi_n_166 = ~(csa_tree_mul_77_11_groupi_n_12 | ((csa_tree_mul_77_11_groupi_n_46
    & n_1321) | (n_1320 & n_1313)));
 assign csa_tree_mul_77_11_groupi_n_165 = ~csa_tree_mul_77_11_groupi_n_104;
 assign csa_tree_mul_77_11_groupi_n_163 = ~csa_tree_mul_77_11_groupi_n_164;
 assign csa_tree_mul_77_11_groupi_n_161 = ~csa_tree_mul_77_11_groupi_n_162;
 assign csa_tree_mul_77_11_groupi_n_160 = ~(csa_tree_mul_77_11_groupi_n_106 | csa_tree_mul_77_11_groupi_n_29);
 assign csa_tree_mul_77_11_groupi_n_159 = ~(csa_tree_mul_77_11_groupi_n_103 | csa_tree_mul_77_11_groupi_n_29);
 assign csa_tree_mul_77_11_groupi_n_158 = ~(csa_tree_mul_77_11_groupi_n_0 | csa_tree_mul_77_11_groupi_n_29);
 assign csa_tree_mul_77_11_groupi_n_164 = ~(csa_tree_mul_77_11_groupi_n_0 & n_1314);
 assign csa_tree_mul_77_11_groupi_n_162 = ~(csa_tree_mul_77_11_groupi_n_105 | csa_tree_mul_77_11_groupi_n_101);
 assign csa_tree_mul_77_11_groupi_n_157 = ~csa_tree_mul_77_11_groupi_n_156;
 assign csa_tree_mul_77_11_groupi_n_155 = ~csa_tree_mul_77_11_groupi_n_154;
 assign csa_tree_mul_77_11_groupi_n_152 = ~csa_tree_mul_77_11_groupi_n_153;
 assign csa_tree_mul_77_11_groupi_n_151 = ~(csa_tree_mul_77_11_groupi_n_105 & csa_tree_mul_77_11_groupi_n_125);
 assign csa_tree_mul_77_11_groupi_n_150 = ~(csa_tree_mul_77_11_groupi_n_56 & ~csa_tree_mul_77_11_groupi_n_106);
 assign csa_tree_mul_77_11_groupi_n_156 = ~(csa_tree_mul_77_11_groupi_n_102 & n_1317);
 assign csa_tree_mul_77_11_groupi_n_154 = ~(csa_tree_mul_77_11_groupi_n_105 & n_1319);
 assign csa_tree_mul_77_11_groupi_n_153 = (csa_tree_mul_77_11_groupi_n_102 | csa_tree_mul_77_11_groupi_n_100);
 assign csa_tree_mul_77_11_groupi_n_143 = ~csa_tree_mul_77_11_groupi_n_142;
 assign csa_tree_mul_77_11_groupi_n_137 = ~csa_tree_mul_77_11_groupi_n_136;
 assign csa_tree_mul_77_11_groupi_n_126 = ~csa_tree_mul_77_11_groupi_n_125;
 assign csa_tree_mul_77_11_groupi_n_119 = ~csa_tree_mul_77_11_groupi_n_118;
 assign csa_tree_mul_77_11_groupi_n_111 = ~csa_tree_mul_77_11_groupi_n_110;
 assign csa_tree_mul_77_11_groupi_n_109 = ~n_1490;
 assign csa_tree_mul_77_11_groupi_n_107 = ~csa_tree_mul_77_11_groupi_n_0;
 assign csa_tree_mul_77_11_groupi_n_105 = ~csa_tree_mul_77_11_groupi_n_106;
 assign csa_tree_mul_77_11_groupi_n_102 = ~csa_tree_mul_77_11_groupi_n_103;
 assign csa_tree_mul_77_11_groupi_n_101 = ~(n_1319 ^ n_1320);
 assign csa_tree_mul_77_11_groupi_n_100 = ~(n_1317 ^ n_1318);
 assign csa_tree_mul_77_11_groupi_n_99 = ~((csa_tree_mul_77_11_groupi_n_26 & n_1315) | (csa_tree_mul_77_11_groupi_n_28
    & n_1316));
 assign csa_tree_mul_77_11_groupi_n_149 = ~((csa_tree_mul_77_11_groupi_n_27 & n_1304) | (csa_tree_mul_77_11_groupi_n_25
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_148 = ~((csa_tree_mul_77_11_groupi_n_12 & n_1311) | (csa_tree_mul_77_11_groupi_n_37
    & n_1319));
 assign csa_tree_mul_77_11_groupi_n_147 = ~((csa_tree_mul_77_11_groupi_n_12 & n_1297) | (csa_tree_mul_77_11_groupi_n_35
    & n_1319));
 assign csa_tree_mul_77_11_groupi_n_98 = ~(n_1350 | csa_tree_mul_77_11_groupi_n_13);
 assign csa_tree_mul_77_11_groupi_n_146 = ~((csa_tree_mul_77_11_groupi_n_27 & n_1310) | (csa_tree_mul_77_11_groupi_n_23
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_145 = ~((csa_tree_mul_77_11_groupi_n_12 & ~n_1309) | (n_1319 & n_1309));
 assign csa_tree_mul_77_11_groupi_n_144 = ~((n_1317 & ~n_1309) | (csa_tree_mul_77_11_groupi_n_27 & n_1309));
 assign csa_tree_mul_77_11_groupi_n_142 = ~((csa_tree_mul_77_11_groupi_n_12 & n_1302) | (csa_tree_mul_77_11_groupi_n_18
    & n_1319));
 assign csa_tree_mul_77_11_groupi_n_141 = ~((csa_tree_mul_77_11_groupi_n_27 & n_1306) | (csa_tree_mul_77_11_groupi_n_16
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_140 = ~((csa_tree_mul_77_11_groupi_n_12 & n_1296) | (csa_tree_mul_77_11_groupi_n_31
    & n_1319));
 assign csa_tree_mul_77_11_groupi_n_139 = ~((csa_tree_mul_77_11_groupi_n_27 & n_1301) | (csa_tree_mul_77_11_groupi_n_34
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_138 = ~((csa_tree_mul_77_11_groupi_n_27 & n_1311) | (csa_tree_mul_77_11_groupi_n_37
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_136 = ~((csa_tree_mul_77_11_groupi_n_27 & ~n_1501) | (n_1317 & n_1501));
 assign csa_tree_mul_77_11_groupi_n_135 = ~((n_1319 & ~n_1502) | (csa_tree_mul_77_11_groupi_n_12 & n_1502));
 assign csa_tree_mul_77_11_groupi_n_134 = ~((csa_tree_mul_77_11_groupi_n_20 & ~csa_tree_mul_77_11_groupi_n_27)
    | (n_1502 & csa_tree_mul_77_11_groupi_n_27));
 assign csa_tree_mul_77_11_groupi_n_133 = ~((csa_tree_mul_77_11_groupi_n_12 & n_1312) | (csa_tree_mul_77_11_groupi_n_22
    & n_1319));
 assign csa_tree_mul_77_11_groupi_n_132 = ~((csa_tree_mul_77_11_groupi_n_27 & n_1297) | (csa_tree_mul_77_11_groupi_n_35
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_131 = ~((csa_tree_mul_77_11_groupi_n_12 & ~n_1501) | (n_1319 & n_1501));
 assign csa_tree_mul_77_11_groupi_n_130 = ~((csa_tree_mul_77_11_groupi_n_27 & n_1299) | (csa_tree_mul_77_11_groupi_n_24
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_129 = ~((csa_tree_mul_77_11_groupi_n_27 & n_1312) | (csa_tree_mul_77_11_groupi_n_22
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_128 = ~((csa_tree_mul_77_11_groupi_n_12 & ~n_1306) | (n_1319 & n_1306));
 assign csa_tree_mul_77_11_groupi_n_127 = ~((csa_tree_mul_77_11_groupi_n_12 & n_1310) | (csa_tree_mul_77_11_groupi_n_23
    & n_1319));
 assign csa_tree_mul_77_11_groupi_n_125 = ~((csa_tree_mul_77_11_groupi_n_12 & ~n_1301) | (n_1319 & n_1301));
 assign csa_tree_mul_77_11_groupi_n_124 = ~((csa_tree_mul_77_11_groupi_n_27 & n_1303) | (csa_tree_mul_77_11_groupi_n_36
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_123 = ~((csa_tree_mul_77_11_groupi_n_12 & n_1299) | (csa_tree_mul_77_11_groupi_n_24
    & n_1319));
 assign csa_tree_mul_77_11_groupi_n_122 = ~((n_1319 | csa_tree_mul_77_11_groupi_n_30) & (n_1294 | csa_tree_mul_77_11_groupi_n_12));
 assign csa_tree_mul_77_11_groupi_n_121 = ~((csa_tree_mul_77_11_groupi_n_12 & n_1300) | (csa_tree_mul_77_11_groupi_n_15
    & n_1319));
 assign csa_tree_mul_77_11_groupi_n_120 = ~((csa_tree_mul_77_11_groupi_n_27 & n_1500) | (csa_tree_mul_77_11_groupi_n_21
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_118 = ~((csa_tree_mul_77_11_groupi_n_12 & n_1295) | (csa_tree_mul_77_11_groupi_n_17
    & n_1319));
 assign csa_tree_mul_77_11_groupi_n_117 = ~((n_1317 | csa_tree_mul_77_11_groupi_n_30) & (n_1294 | csa_tree_mul_77_11_groupi_n_27));
 assign csa_tree_mul_77_11_groupi_n_116 = ~((csa_tree_mul_77_11_groupi_n_27 & n_1298) | (csa_tree_mul_77_11_groupi_n_32
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_115 = ~((csa_tree_mul_77_11_groupi_n_27 & n_1296) | (csa_tree_mul_77_11_groupi_n_31
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_114 = ~((csa_tree_mul_77_11_groupi_n_12 & n_1298) | (csa_tree_mul_77_11_groupi_n_32
    & n_1319));
 assign csa_tree_mul_77_11_groupi_n_113 = ~((csa_tree_mul_77_11_groupi_n_12 & n_1303) | (csa_tree_mul_77_11_groupi_n_36
    & n_1319));
 assign csa_tree_mul_77_11_groupi_n_112 = ~((csa_tree_mul_77_11_groupi_n_27 & n_1302) | (csa_tree_mul_77_11_groupi_n_18
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_110 = ~((csa_tree_mul_77_11_groupi_n_27 & n_1295) | (csa_tree_mul_77_11_groupi_n_17
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_106 = ((n_1320 | csa_tree_mul_77_11_groupi_n_13) & (n_1321 | csa_tree_mul_77_11_groupi_n_38));
 assign csa_tree_mul_77_11_groupi_n_104 = ~(n_1317 ^ n_1316);
 assign csa_tree_mul_77_11_groupi_n_103 = ~(n_1318 ^ n_1319);
 assign csa_tree_mul_77_11_groupi_n_90 = ~csa_tree_mul_77_11_groupi_n_89;
 assign csa_tree_mul_77_11_groupi_n_83 = ~csa_tree_mul_77_11_groupi_n_82;
 assign csa_tree_mul_77_11_groupi_n_75 = ~csa_tree_mul_77_11_groupi_n_74;
 assign csa_tree_mul_77_11_groupi_n_60 = ~csa_tree_mul_77_11_groupi_n_59;
 assign csa_tree_mul_77_11_groupi_n_57 = ~csa_tree_mul_77_11_groupi_n_56;
 assign csa_tree_mul_77_11_groupi_n_52 = ~((csa_tree_mul_77_11_groupi_n_13 & n_1313) | (csa_tree_mul_77_11_groupi_n_29
    & n_1321));
 assign csa_tree_mul_77_11_groupi_n_51 = ~((csa_tree_mul_77_11_groupi_n_12 & n_1313) | (csa_tree_mul_77_11_groupi_n_29
    & n_1319));
 assign csa_tree_mul_77_11_groupi_n_50 = ~((csa_tree_mul_77_11_groupi_n_27 & n_1313) | (csa_tree_mul_77_11_groupi_n_29
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_49 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1313) | (csa_tree_mul_77_11_groupi_n_29
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_97 = ~((n_1321 & ~n_1304) | (csa_tree_mul_77_11_groupi_n_13 & n_1304));
 assign csa_tree_mul_77_11_groupi_n_96 = ~((csa_tree_mul_77_11_groupi_n_13 & n_1312) | (csa_tree_mul_77_11_groupi_n_22
    & n_1321));
 assign csa_tree_mul_77_11_groupi_n_95 = ~((n_1321 & ~n_1309) | (csa_tree_mul_77_11_groupi_n_13 & n_1309));
 assign csa_tree_mul_77_11_groupi_n_94 = ~((csa_tree_mul_77_11_groupi_n_13 & n_1297) | (csa_tree_mul_77_11_groupi_n_35
    & n_1321));
 assign csa_tree_mul_77_11_groupi_n_93 = ~((n_1321 & ~n_1298) | (csa_tree_mul_77_11_groupi_n_13 & n_1298));
 assign csa_tree_mul_77_11_groupi_n_92 = ~((n_1321 & ~n_1501) | (csa_tree_mul_77_11_groupi_n_13 & n_1501));
 assign csa_tree_mul_77_11_groupi_n_91 = ~((csa_tree_mul_77_11_groupi_n_13 & n_1295) | (csa_tree_mul_77_11_groupi_n_17
    & n_1321));
 assign csa_tree_mul_77_11_groupi_n_89 = ~((csa_tree_mul_77_11_groupi_n_13 & n_1294) | (csa_tree_mul_77_11_groupi_n_30
    & n_1321));
 assign csa_tree_mul_77_11_groupi_n_88 = ~((csa_tree_mul_77_11_groupi_n_15 & ~csa_tree_mul_77_11_groupi_n_13)
    | (n_1300 & csa_tree_mul_77_11_groupi_n_13));
 assign csa_tree_mul_77_11_groupi_n_87 = ~((n_1321 & ~n_1301) | (csa_tree_mul_77_11_groupi_n_13 & n_1301));
 assign csa_tree_mul_77_11_groupi_n_86 = ~((csa_tree_mul_77_11_groupi_n_13 & n_1296) | (csa_tree_mul_77_11_groupi_n_31
    & n_1321));
 assign csa_tree_mul_77_11_groupi_n_85 = ~((csa_tree_mul_77_11_groupi_n_13 & n_1311) | (csa_tree_mul_77_11_groupi_n_37
    & n_1321));
 assign csa_tree_mul_77_11_groupi_n_84 = ~((n_1321 & ~n_1502) | (csa_tree_mul_77_11_groupi_n_13 & n_1502));
 assign csa_tree_mul_77_11_groupi_n_82 = ~((csa_tree_mul_77_11_groupi_n_13 & ~n_1303) | (n_1321 & n_1303));
 assign csa_tree_mul_77_11_groupi_n_81 = ~((csa_tree_mul_77_11_groupi_n_13 & n_1310) | (csa_tree_mul_77_11_groupi_n_23
    & n_1321));
 assign csa_tree_mul_77_11_groupi_n_80 = ~((n_1321 & ~n_1500) | (csa_tree_mul_77_11_groupi_n_13 & n_1500));
 assign csa_tree_mul_77_11_groupi_n_79 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1297) | (csa_tree_mul_77_11_groupi_n_35
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_78 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1306) | (csa_tree_mul_77_11_groupi_n_16
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_77 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1296) | (csa_tree_mul_77_11_groupi_n_31
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_76 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1303) | (csa_tree_mul_77_11_groupi_n_36
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_74 = ~((csa_tree_mul_77_11_groupi_n_28 & ~n_1309) | (n_1315 & n_1309));
 assign csa_tree_mul_77_11_groupi_n_73 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1311) | (csa_tree_mul_77_11_groupi_n_37
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_72 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1300) | (csa_tree_mul_77_11_groupi_n_15
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_71 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1310) | (csa_tree_mul_77_11_groupi_n_23
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_70 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1299) | (csa_tree_mul_77_11_groupi_n_24
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_69 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1500) | (csa_tree_mul_77_11_groupi_n_21
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_68 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1302) | (csa_tree_mul_77_11_groupi_n_18
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_67 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1304) | (csa_tree_mul_77_11_groupi_n_25
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_66 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1312) | (csa_tree_mul_77_11_groupi_n_22
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_65 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1301) | (csa_tree_mul_77_11_groupi_n_34
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_64 = ~((n_1315 | csa_tree_mul_77_11_groupi_n_30) & (n_1294 | csa_tree_mul_77_11_groupi_n_28));
 assign csa_tree_mul_77_11_groupi_n_63 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1298) | (csa_tree_mul_77_11_groupi_n_32
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_62 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1501) | (csa_tree_mul_77_11_groupi_n_33
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_61 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1502) | (csa_tree_mul_77_11_groupi_n_20
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_59 = ~((csa_tree_mul_77_11_groupi_n_28 & n_1295) | (csa_tree_mul_77_11_groupi_n_17
    & n_1315));
 assign csa_tree_mul_77_11_groupi_n_58 = ~((csa_tree_mul_77_11_groupi_n_27 & n_1300) | (csa_tree_mul_77_11_groupi_n_15
    & n_1317));
 assign csa_tree_mul_77_11_groupi_n_56 = ~((csa_tree_mul_77_11_groupi_n_12 & ~n_1304) | (n_1319 & n_1304));
 assign csa_tree_mul_77_11_groupi_n_55 = ~((n_1321 & ~n_1302) | (csa_tree_mul_77_11_groupi_n_13 & n_1302));
 assign csa_tree_mul_77_11_groupi_n_54 = ~((csa_tree_mul_77_11_groupi_n_13 & n_1299) | (csa_tree_mul_77_11_groupi_n_24
    & n_1321));
 assign csa_tree_mul_77_11_groupi_n_47 = ~(csa_tree_mul_77_11_groupi_n_27 & csa_tree_mul_77_11_groupi_n_26);
 assign csa_tree_mul_77_11_groupi_n_46 = ~(csa_tree_mul_77_11_groupi_n_38 & csa_tree_mul_77_11_groupi_n_29);
 assign n_1350 = (n_1322 & n_1313);
 assign csa_tree_mul_77_11_groupi_n_40 = ~(csa_tree_mul_77_11_groupi_n_12 & csa_tree_mul_77_11_groupi_n_29);
 assign csa_tree_mul_77_11_groupi_n_39 = ~(n_1322 & n_1321);
 assign csa_tree_mul_77_11_groupi_n_38 = ~n_1320;
 assign csa_tree_mul_77_11_groupi_n_37 = ~n_1311;
 assign csa_tree_mul_77_11_groupi_n_36 = ~n_1303;
 assign csa_tree_mul_77_11_groupi_n_35 = ~n_1297;
 assign csa_tree_mul_77_11_groupi_n_34 = ~n_1301;
 assign csa_tree_mul_77_11_groupi_n_33 = ~n_1501;
 assign csa_tree_mul_77_11_groupi_n_32 = ~n_1298;
 assign csa_tree_mul_77_11_groupi_n_31 = ~n_1296;
 assign csa_tree_mul_77_11_groupi_n_30 = ~n_1294;
 assign csa_tree_mul_77_11_groupi_n_29 = ~n_1313;
 assign csa_tree_mul_77_11_groupi_n_28 = ~n_1315;
 assign csa_tree_mul_77_11_groupi_n_27 = ~n_1317;
 assign csa_tree_mul_77_11_groupi_n_26 = ~n_1316;
 assign csa_tree_mul_77_11_groupi_n_25 = ~n_1304;
 assign csa_tree_mul_77_11_groupi_n_24 = ~n_1299;
 assign csa_tree_mul_77_11_groupi_n_23 = ~n_1310;
 assign csa_tree_mul_77_11_groupi_n_22 = ~n_1312;
 assign csa_tree_mul_77_11_groupi_n_21 = ~n_1500;
 assign csa_tree_mul_77_11_groupi_n_20 = ~n_1502;
 assign csa_tree_mul_77_11_groupi_n_19 = ~n_1309;
 assign csa_tree_mul_77_11_groupi_n_18 = ~n_1302;
 assign csa_tree_mul_77_11_groupi_n_17 = ~n_1295;
 assign csa_tree_mul_77_11_groupi_n_16 = ~n_1306;
 assign csa_tree_mul_77_11_groupi_n_15 = ~n_1300;
 assign csa_tree_mul_77_11_groupi_n_14 = ~n_1322;
 assign csa_tree_mul_77_11_groupi_n_13 = ~n_1321;
 assign csa_tree_mul_77_11_groupi_n_12 = ~n_1319;
 assign csa_tree_mul_77_11_groupi_n_9 = (csa_tree_mul_77_11_groupi_n_500 | csa_tree_mul_77_11_groupi_n_7);
 assign csa_tree_mul_77_11_groupi_n_7 = (csa_tree_mul_77_11_groupi_n_478 & csa_tree_mul_77_11_groupi_n_454);
 assign csa_tree_mul_77_11_groupi_n_6 = ~(csa_tree_mul_77_11_groupi_n_462 | ~csa_tree_mul_77_11_groupi_n_461);
 assign csa_tree_mul_77_11_groupi_n_5 = ~(csa_tree_mul_77_11_groupi_n_3 & ~csa_tree_mul_77_11_groupi_n_442);
 assign csa_tree_mul_77_11_groupi_n_3 = ~(csa_tree_mul_77_11_groupi_n_444 & ~csa_tree_mul_77_11_groupi_n_385);
 assign csa_tree_mul_77_11_groupi_n_2 = ~(csa_tree_mul_77_11_groupi_n_295 ^ csa_tree_mul_77_11_groupi_n_365);
 assign csa_tree_mul_77_11_groupi_n_1 = (csa_tree_mul_77_11_groupi_n_92 | n_1489);
 assign csa_tree_mul_77_11_groupi_n_0 = ((csa_tree_mul_77_11_groupi_n_28 & ~n_1314) | (n_1315 & n_1314));
 assign final_adder_add_69_2_n_12 = ((final_adder_add_69_2_n_10 & {in1[6]}) | (({in1[6]} & {in2[6]})
    | ({in2[6]} & final_adder_add_69_2_n_10)));
 assign n_1432 = ({in1[6]} ^ ({in2[6]} ^ final_adder_add_69_2_n_10));
 assign final_adder_add_69_2_n_8 = ((final_adder_add_69_2_n_6 & {in1[4]}) | (({in1[4]} & {in2[4]}) |
    ({in2[4]} & final_adder_add_69_2_n_6)));
 assign n_1434 = ({in1[4]} ^ ({in2[4]} ^ final_adder_add_69_2_n_6));
 assign final_adder_add_69_2_n_4 = ((final_adder_add_69_2_n_2 & {in1[2]}) | (({in1[2]} & {in2[2]}) |
    ({in2[2]} & final_adder_add_69_2_n_2)));
 assign n_1436 = ({in1[2]} ^ ({in2[2]} ^ final_adder_add_69_2_n_2));
 assign final_adder_add_86_2_n_49 = ((final_adder_add_86_2_n_47 & n_1355) | ((n_1355 & n_1386) | (n_1386
    & final_adder_add_86_2_n_47)));
 assign n_1411 = (n_1355 ^ (n_1386 ^ final_adder_add_86_2_n_47));
 assign final_adder_add_86_2_n_47 = ((final_adder_add_86_2_n_45 & n_1356) | ((n_1356 & n_1387) | (n_1387
    & final_adder_add_86_2_n_45)));
 assign n_1412 = (n_1356 ^ (n_1387 ^ final_adder_add_86_2_n_45));
 assign final_adder_add_86_2_n_45 = ((final_adder_add_86_2_n_43 & n_1357) | ((n_1357 & n_1388) | (n_1388
    & final_adder_add_86_2_n_43)));
 assign n_1413 = (n_1357 ^ (n_1388 ^ final_adder_add_86_2_n_43));
 assign final_adder_add_86_2_n_43 = ((final_adder_add_86_2_n_41 & n_1358) | ((n_1358 & n_1389) | (n_1389
    & final_adder_add_86_2_n_41)));
 assign n_1414 = (n_1358 ^ (n_1389 ^ final_adder_add_86_2_n_41));
 assign final_adder_add_86_2_n_41 = ((final_adder_add_86_2_n_39 & n_1359) | ((n_1359 & n_1390) | (n_1390
    & final_adder_add_86_2_n_39)));
 assign n_1415 = (n_1359 ^ (n_1390 ^ final_adder_add_86_2_n_39));
 assign final_adder_add_86_2_n_39 = ((final_adder_add_86_2_n_37 & n_1360) | ((n_1360 & n_1391) | (n_1391
    & final_adder_add_86_2_n_37)));
 assign n_1416 = (n_1360 ^ (n_1391 ^ final_adder_add_86_2_n_37));
 assign final_adder_add_86_2_n_37 = ((final_adder_add_86_2_n_35 & n_1392) | ((n_1392 & n_1361) | (n_1361
    & final_adder_add_86_2_n_35)));
 assign n_1417 = (n_1392 ^ (n_1361 ^ final_adder_add_86_2_n_35));
 assign final_adder_add_86_2_n_35 = ((final_adder_add_86_2_n_33 & n_1362) | ((n_1362 & n_1393) | (n_1393
    & final_adder_add_86_2_n_33)));
 assign n_1418 = (n_1362 ^ (n_1393 ^ final_adder_add_86_2_n_33));
 assign final_adder_add_86_2_n_33 = ((final_adder_add_86_2_n_31 & n_1363) | ((n_1363 & n_1394) | (n_1394
    & final_adder_add_86_2_n_31)));
 assign n_1419 = (n_1363 ^ (n_1394 ^ final_adder_add_86_2_n_31));
 assign final_adder_add_86_2_n_31 = ((final_adder_add_86_2_n_29 & n_1364) | ((n_1364 & n_1395) | (n_1395
    & final_adder_add_86_2_n_29)));
 assign n_1420 = (n_1364 ^ (n_1395 ^ final_adder_add_86_2_n_29));
 assign final_adder_add_86_2_n_29 = ((final_adder_add_86_2_n_27 & n_1365) | ((n_1365 & n_1396) | (n_1396
    & final_adder_add_86_2_n_27)));
 assign n_1421 = (n_1365 ^ (n_1396 ^ final_adder_add_86_2_n_27));
 assign final_adder_add_86_2_n_27 = ((final_adder_add_86_2_n_25 & n_1366) | ((n_1366 & n_1397) | (n_1397
    & final_adder_add_86_2_n_25)));
 assign n_1422 = (n_1366 ^ (n_1397 ^ final_adder_add_86_2_n_25));
 assign final_adder_add_86_2_n_25 = ((final_adder_add_86_2_n_23 & n_1367) | ((n_1367 & n_1398) | (n_1398
    & final_adder_add_86_2_n_23)));
 assign n_1423 = (n_1367 ^ (n_1398 ^ final_adder_add_86_2_n_23));
 assign final_adder_add_86_2_n_23 = ((final_adder_add_86_2_n_21 & n_1368) | ((n_1368 & n_1399) | (n_1399
    & final_adder_add_86_2_n_21)));
 assign n_1424 = (n_1368 ^ (n_1399 ^ final_adder_add_86_2_n_21));
 assign final_adder_add_86_2_n_21 = ((final_adder_add_86_2_n_19 & n_1369) | ((n_1369 & n_1400) | (n_1400
    & final_adder_add_86_2_n_19)));
 assign n_1425 = (n_1369 ^ (n_1400 ^ final_adder_add_86_2_n_19));
 assign final_adder_add_86_2_n_3 = ((final_adder_add_86_2_n_1 & n_1376) | ((n_1376 & n_1406) | (n_1406
    & final_adder_add_86_2_n_1)));
 assign n_1428 = (n_1376 ^ (n_1406 ^ final_adder_add_86_2_n_1));
 assign final_adder_add_86_2_n_1 = (n_1407 & n_1377);
 assign n_1429 = (n_1407 ^ n_1377);
 assign n_446 = ((csa_tree_add_92_2_groupi_n_93 & n_448) | ((n_448 & n_674) | (n_674 & csa_tree_add_92_2_groupi_n_93)));
 assign n_445 = (n_448 ^ (n_674 ^ csa_tree_add_92_2_groupi_n_93));
 assign n_448 = ((csa_tree_add_92_2_groupi_n_94 & n_450) | ((n_450 & csa_tree_add_92_2_groupi_n_79) |
    (csa_tree_add_92_2_groupi_n_79 & csa_tree_add_92_2_groupi_n_94)));
 assign n_447 = (n_450 ^ (csa_tree_add_92_2_groupi_n_79 ^ csa_tree_add_92_2_groupi_n_94));
 assign n_454 = ((n_1012 & n_459) | ((n_459 & csa_tree_add_106_2_groupi_n_1081) | (csa_tree_add_106_2_groupi_n_1081
    & n_1012)));
 assign n_453 = (n_459 ^ (csa_tree_add_106_2_groupi_n_1081 ^ n_1012));
 assign n_450 = ((csa_tree_add_92_2_groupi_n_80 & n_452) | ((n_452 & csa_tree_add_92_2_groupi_n_83) |
    (csa_tree_add_92_2_groupi_n_83 & csa_tree_add_92_2_groupi_n_80)));
 assign n_449 = (n_452 ^ (csa_tree_add_92_2_groupi_n_83 ^ csa_tree_add_92_2_groupi_n_80));
 assign n_457 = ~((n_458 & n_465) | (n_1143 & stall));
 assign n_459 = ((n_463 & csa_tree_add_106_2_groupi_n_1082) | ((csa_tree_add_106_2_groupi_n_1082 & csa_tree_add_106_2_groupi_n_1051)
    | (csa_tree_add_106_2_groupi_n_1051 & n_463)));
 assign n_458 = (csa_tree_add_106_2_groupi_n_1082 ^ (csa_tree_add_106_2_groupi_n_1051 ^ n_463));
 assign n_452 = ((csa_tree_add_92_2_groupi_n_87 & n_456) | ((n_456 & csa_tree_add_92_2_groupi_n_84) |
    (csa_tree_add_92_2_groupi_n_84 & csa_tree_add_92_2_groupi_n_87)));
 assign n_451 = (n_456 ^ (csa_tree_add_92_2_groupi_n_84 ^ csa_tree_add_92_2_groupi_n_87));
 assign n_463 = ((n_467 & csa_tree_add_106_2_groupi_n_1052) | ((csa_tree_add_106_2_groupi_n_1052 & csa_tree_add_106_2_groupi_n_1114)
    | (csa_tree_add_106_2_groupi_n_1114 & n_467)));
 assign n_462 = (csa_tree_add_106_2_groupi_n_1052 ^ (csa_tree_add_106_2_groupi_n_1114 ^ n_467));
 assign n_456 = ((csa_tree_add_92_2_groupi_n_88 & n_461) | ((n_461 & csa_tree_add_92_2_groupi_n_67) |
    (csa_tree_add_92_2_groupi_n_67 & csa_tree_add_92_2_groupi_n_88)));
 assign n_455 = (n_461 ^ (csa_tree_add_92_2_groupi_n_67 ^ csa_tree_add_92_2_groupi_n_88));
 assign n_464 = ~((n_466 & n_465) | (n_1146 & stall));
 assign n_467 = ((n_471 & csa_tree_add_106_2_groupi_n_1115) | ((csa_tree_add_106_2_groupi_n_1115 & csa_tree_add_106_2_groupi_n_1108)
    | (csa_tree_add_106_2_groupi_n_1108 & n_471)));
 assign n_466 = (csa_tree_add_106_2_groupi_n_1115 ^ (csa_tree_add_106_2_groupi_n_1108 ^ n_471));
 assign n_461 = ((csa_tree_add_92_2_groupi_n_68 & n_469) | ((n_469 & csa_tree_add_92_2_groupi_n_85) |
    (csa_tree_add_92_2_groupi_n_85 & csa_tree_add_92_2_groupi_n_68)));
 assign n_460 = (n_469 ^ (csa_tree_add_92_2_groupi_n_85 ^ csa_tree_add_92_2_groupi_n_68));
 assign n_471 = ((n_475 & csa_tree_add_106_2_groupi_n_1109) | ((csa_tree_add_106_2_groupi_n_1109 & csa_tree_add_106_2_groupi_n_1110)
    | (csa_tree_add_106_2_groupi_n_1110 & n_475)));
 assign n_470 = (csa_tree_add_106_2_groupi_n_1109 ^ (csa_tree_add_106_2_groupi_n_1110 ^ n_475));
 assign n_469 = ((csa_tree_add_92_2_groupi_n_86 & n_473) | ((n_473 & csa_tree_add_92_2_groupi_n_71) |
    (csa_tree_add_92_2_groupi_n_71 & csa_tree_add_92_2_groupi_n_86)));
 assign n_468 = (n_473 ^ (csa_tree_add_92_2_groupi_n_71 ^ csa_tree_add_92_2_groupi_n_86));
 assign n_475 = ((n_477 & csa_tree_add_106_2_groupi_n_1111) | ((csa_tree_add_106_2_groupi_n_1111 & csa_tree_add_106_2_groupi_n_1120)
    | (csa_tree_add_106_2_groupi_n_1120 & n_477)));
 assign n_474 = (csa_tree_add_106_2_groupi_n_1111 ^ (csa_tree_add_106_2_groupi_n_1120 ^ n_477));
 assign n_473 = ((csa_tree_add_92_2_groupi_n_73 & n_479) | ((n_479 & csa_tree_add_92_2_groupi_n_72) |
    (csa_tree_add_92_2_groupi_n_72 & csa_tree_add_92_2_groupi_n_73)));
 assign n_472 = (n_479 ^ (csa_tree_add_92_2_groupi_n_72 ^ csa_tree_add_92_2_groupi_n_73));
 assign n_477 = ((n_481 & csa_tree_add_106_2_groupi_n_1121) | ((csa_tree_add_106_2_groupi_n_1121 & csa_tree_add_106_2_groupi_n_1118)
    | (csa_tree_add_106_2_groupi_n_1118 & n_481)));
 assign n_476 = (csa_tree_add_106_2_groupi_n_1121 ^ (csa_tree_add_106_2_groupi_n_1118 ^ n_481));
 assign n_479 = ((csa_tree_add_92_2_groupi_n_74 & n_483) | ((n_483 & csa_tree_add_92_2_groupi_n_69) |
    (csa_tree_add_92_2_groupi_n_69 & csa_tree_add_92_2_groupi_n_74)));
 assign n_478 = (n_483 ^ (csa_tree_add_92_2_groupi_n_69 ^ csa_tree_add_92_2_groupi_n_74));
 assign n_481 = ((n_485 & csa_tree_add_106_2_groupi_n_1119) | ((csa_tree_add_106_2_groupi_n_1119 & csa_tree_add_106_2_groupi_n_1112)
    | (csa_tree_add_106_2_groupi_n_1112 & n_485)));
 assign n_480 = (csa_tree_add_106_2_groupi_n_1119 ^ (csa_tree_add_106_2_groupi_n_1112 ^ n_485));
 assign n_483 = ((csa_tree_add_92_2_groupi_n_70 & n_487) | ((n_487 & csa_tree_add_92_2_groupi_n_77) |
    (csa_tree_add_92_2_groupi_n_77 & csa_tree_add_92_2_groupi_n_70)));
 assign n_482 = (n_487 ^ (csa_tree_add_92_2_groupi_n_77 ^ csa_tree_add_92_2_groupi_n_70));
 assign n_485 = ((csa_tree_add_106_2_groupi_n_1113 & n_489) | ((n_489 & csa_tree_add_106_2_groupi_n_1106)
    | (csa_tree_add_106_2_groupi_n_1106 & csa_tree_add_106_2_groupi_n_1113)));
 assign n_484 = (n_489 ^ (csa_tree_add_106_2_groupi_n_1106 ^ csa_tree_add_106_2_groupi_n_1113));
 assign n_487 = ((csa_tree_add_92_2_groupi_n_176 & n_491) | ((n_491 & csa_tree_add_92_2_groupi_n_78)
    | (csa_tree_add_92_2_groupi_n_78 & csa_tree_add_92_2_groupi_n_176)));
 assign n_486 = (n_491 ^ (csa_tree_add_92_2_groupi_n_78 ^ csa_tree_add_92_2_groupi_n_176));
 assign n_489 = ((csa_tree_add_106_2_groupi_n_1107 & n_493) | ((n_493 & csa_tree_add_106_2_groupi_n_1098)
    | (csa_tree_add_106_2_groupi_n_1098 & csa_tree_add_106_2_groupi_n_1107)));
 assign n_488 = (n_493 ^ (csa_tree_add_106_2_groupi_n_1098 ^ csa_tree_add_106_2_groupi_n_1107));
 assign n_491 = ((csa_tree_add_92_2_groupi_n_177 & n_498) | ((n_498 & csa_tree_add_92_2_groupi_n_204)
    | (csa_tree_add_92_2_groupi_n_204 & csa_tree_add_92_2_groupi_n_177)));
 assign n_490 = (n_498 ^ (csa_tree_add_92_2_groupi_n_204 ^ csa_tree_add_92_2_groupi_n_177));
 assign n_493 = ((n_496 & csa_tree_add_106_2_groupi_n_1099) | ((csa_tree_add_106_2_groupi_n_1099 & csa_tree_add_106_2_groupi_n_1094)
    | (csa_tree_add_106_2_groupi_n_1094 & n_496)));
 assign n_492 = (csa_tree_add_106_2_groupi_n_1099 ^ (csa_tree_add_106_2_groupi_n_1094 ^ n_496));
 assign n_498 = ((n_505 & csa_tree_add_92_2_groupi_n_205) | ((csa_tree_add_92_2_groupi_n_205 & csa_tree_add_92_2_groupi_n_210)
    | (csa_tree_add_92_2_groupi_n_210 & n_505)));
 assign n_497 = (csa_tree_add_92_2_groupi_n_205 ^ (csa_tree_add_92_2_groupi_n_210 ^ n_505));
 assign n_494 = ~((n_495 & n_465) | (n_201 & stall));
 assign n_496 = ((n_502 & csa_tree_add_106_2_groupi_n_1095) | ((csa_tree_add_106_2_groupi_n_1095 & csa_tree_add_106_2_groupi_n_1063)
    | (csa_tree_add_106_2_groupi_n_1063 & n_502)));
 assign n_495 = (csa_tree_add_106_2_groupi_n_1095 ^ (csa_tree_add_106_2_groupi_n_1063 ^ n_502));
 assign n_505 = ((n_512 & csa_tree_add_92_2_groupi_n_211) | ((csa_tree_add_92_2_groupi_n_211 & csa_tree_add_92_2_groupi_n_220)
    | (csa_tree_add_92_2_groupi_n_220 & n_512)));
 assign n_504 = (csa_tree_add_92_2_groupi_n_211 ^ (csa_tree_add_92_2_groupi_n_220 ^ n_512));
 assign n_499 = ~(n_500 ^ n_503);
 assign n_502 = ((n_509 & csa_tree_add_106_2_groupi_n_1064) | ((csa_tree_add_106_2_groupi_n_1064 & csa_tree_add_106_2_groupi_n_1039)
    | (csa_tree_add_106_2_groupi_n_1039 & n_509)));
 assign n_500 = (csa_tree_add_106_2_groupi_n_1064 ^ (csa_tree_add_106_2_groupi_n_1039 ^ n_509));
 assign n_512 = ((n_522 & csa_tree_add_92_2_groupi_n_221) | ((csa_tree_add_92_2_groupi_n_221 & csa_tree_add_92_2_groupi_n_226)
    | (csa_tree_add_92_2_groupi_n_226 & n_522)));
 assign n_511 = (csa_tree_add_92_2_groupi_n_221 ^ (csa_tree_add_92_2_groupi_n_226 ^ n_522));
 assign n_501 = ~((n_506 & n_465) | (n_1157 & stall));
 assign n_509 = ((n_518 & csa_tree_add_106_2_groupi_n_1040) | ((csa_tree_add_106_2_groupi_n_1040 & csa_tree_add_106_2_groupi_n_1008)
    | (csa_tree_add_106_2_groupi_n_1008 & n_518)));
 assign n_503 = (csa_tree_add_106_2_groupi_n_1040 ^ (csa_tree_add_106_2_groupi_n_1008 ^ n_518));
 assign n_507 = ((n_1015 & n_517) | ((n_517 & csa_tree_add_92_2_groupi_n_202) | (csa_tree_add_92_2_groupi_n_202
    & n_1015)));
 assign n_506 = (n_517 ^ (csa_tree_add_92_2_groupi_n_202 ^ n_1015));
 assign n_508 = ~((n_513 & n_465) | (n_800 & stall));
 assign n_522 = ((n_533 & csa_tree_add_92_2_groupi_n_227) | ((csa_tree_add_92_2_groupi_n_227 & n_566)
    | (n_566 & n_533)));
 assign n_521 = (csa_tree_add_92_2_groupi_n_227 ^ (n_566 ^ n_533));
 assign n_513 = ~(n_514 ^ n_520);
 assign n_515 = ~(n_523 ^ n_780);
 assign n_510 = ~((n_516 & n_465) | (n_1158 & stall));
 assign n_518 = ((n_528 & csa_tree_add_106_2_groupi_n_1010) | ((csa_tree_add_106_2_groupi_n_1010 & n_555)
    | (n_555 & n_528)));
 assign n_514 = (csa_tree_add_106_2_groupi_n_1010 ^ (n_555 ^ n_528));
 assign n_519 = ~(n_690 & (n_689 | n_526));
 assign n_523 = ~(n_527 ^ n_1370);
 assign n_517 = ((n_525 & csa_tree_add_92_2_groupi_n_203) | ((csa_tree_add_92_2_groupi_n_203 & csa_tree_add_92_2_groupi_n_192)
    | (csa_tree_add_92_2_groupi_n_192 & n_525)));
 assign n_516 = (csa_tree_add_92_2_groupi_n_203 ^ (csa_tree_add_92_2_groupi_n_192 ^ n_525));
 assign mul_109_11_n_553 = ~(mul_109_11_n_31 | ((n_1456 & n_362) | (mul_109_11_n_64 & n_1455)));
 assign n_526 = ~n_527;
 assign n_530 = ~(n_1016 ^ n_531);
 assign n_527 = ~(n_1156 & ~(n_1155 & n_531));
 assign csa_tree_add_106_2_groupi_n_1085 = ((n_529 & csa_tree_add_106_2_groupi_n_1023) | ((csa_tree_add_106_2_groupi_n_1023
    & n_50) | (n_50 & n_529)));
 assign csa_tree_add_106_2_groupi_n_1086 = (csa_tree_add_106_2_groupi_n_1023 ^ (n_50 ^ n_529));
 assign n_533 = ((n_565 & n_559) | ((n_559 & n_656) | (n_656 & n_565)));
 assign n_532 = (n_559 ^ (n_656 ^ n_565));
 assign n_525 = ((n_537 & csa_tree_add_92_2_groupi_n_193) | ((csa_tree_add_92_2_groupi_n_193 & csa_tree_add_92_2_groupi_n_174)
    | (csa_tree_add_92_2_groupi_n_174 & n_537)));
 assign n_524 = (csa_tree_add_92_2_groupi_n_193 ^ (csa_tree_add_92_2_groupi_n_174 ^ n_537));
 assign n_531 = ((n_561 & n_1402) | ((n_1402 & n_1372) | (n_1372 & n_561)));
 assign n_535 = (n_1402 ^ (n_1372 ^ n_561));
 assign csa_tree_add_106_2_groupi_n_1150 = ((n_974 & n_562) | ((n_562 & n_17) | (n_17 & n_974)));
 assign n_1455 = (n_562 ^ (n_17 ^ n_974));
 assign n_528 = ((n_554 & n_553) | ((n_553 & n_606) | (n_606 & n_554)));
 assign n_520 = (n_553 ^ (n_606 ^ n_554));
 assign csa_tree_add_106_2_groupi_n_962 = ((n_545 & n_543) | ((n_543 & n_48) | (n_48 & n_545)));
 assign csa_tree_add_106_2_groupi_n_963 = (n_543 ^ (n_48 ^ n_545));
 assign csa_tree_add_106_2_groupi_n_972 = ((n_57 & n_534) | ((n_534 & n_53) | (n_53 & n_57)));
 assign csa_tree_add_106_2_groupi_n_973 = (n_534 ^ (n_53 ^ n_57));
 assign n_559 = ((n_655 & n_659) | ((n_659 & n_1147) | (n_1147 & n_655)));
 assign n_558 = (n_659 ^ (n_1147 ^ n_655));
 assign csa_tree_add_106_2_groupi_n_1016 = ((n_54 & n_551) | ((n_551 & n_49) | (n_49 & n_54)));
 assign csa_tree_add_106_2_groupi_n_1017 = (n_551 ^ (n_49 ^ n_54));
 assign n_529 = ((n_610 & n_550) | ((n_550 & n_55) | (n_55 & n_610)));
 assign csa_tree_add_106_2_groupi_n_1027 = (n_550 ^ (n_55 ^ n_610));
 assign mul_109_11_n_101 = ~((n_1456 | n_1) & (mul_109_11_n_28 | n_751));
 assign mul_109_11_n_111 = ~((n_1456 | n_106) & (mul_109_11_n_28 | n_749));
 assign mul_109_11_n_75 = ~((n_1456 | n_362) & (mul_109_11_n_28 | mul_109_11_n_38));
 assign mul_109_11_n_100 = ~((n_1456 | n_433) & (mul_109_11_n_28 | n_777));
 assign mul_109_11_n_92 = ~((n_1456 | n_90) & (mul_109_11_n_28 | n_743));
 assign mul_109_11_n_94 = ~((n_1456 | n_96) & (mul_109_11_n_28 | n_746));
 assign mul_109_11_n_95 = ~((n_1456 | n_95) & (mul_109_11_n_28 | n_745));
 assign mul_109_11_n_93 = ~((n_1456 | n_92) & (mul_109_11_n_28 | n_744));
 assign mul_109_11_n_106 = ~((n_1456 | n_97) & (mul_109_11_n_28 | n_747));
 assign mul_109_11_n_73 = ~((n_1456 | n_748) & (mul_109_11_n_28 | n_98));
 assign n_537 = ((n_568 & csa_tree_add_92_2_groupi_n_175) | ((csa_tree_add_92_2_groupi_n_175 & csa_tree_add_92_2_groupi_n_148)
    | (csa_tree_add_92_2_groupi_n_148 & n_568)));
 assign n_536 = (csa_tree_add_92_2_groupi_n_175 ^ (csa_tree_add_92_2_groupi_n_148 ^ n_568));
 assign n_561 = ((n_1373 & n_1403) | ((n_1403 & n_661) | (n_661 & n_1373)));
 assign n_560 = (n_1403 ^ (n_661 ^ n_1373));
 assign n_553 = ((n_605 & n_602) | ((n_602 & n_133) | (n_133 & n_605)));
 assign n_552 = (n_602 ^ (n_133 ^ n_605));
 assign n_562 = ((n_27 & n_664) | ((n_664 & n_18) | (n_18 & n_27)));
 assign n_1456 = (n_664 ^ (n_18 ^ n_27));
 assign csa_tree_add_106_2_groupi_n_970 = ((n_831 & n_612) | ((n_612 & n_163) | (n_163 & n_831)));
 assign csa_tree_add_106_2_groupi_n_971 = (n_612 ^ (n_163 ^ n_831));
 assign n_539 = ((n_190 & n_580) | ((n_580 & csa_tree_add_106_2_groupi_n_818) | (csa_tree_add_106_2_groupi_n_818
    & n_190)));
 assign n_538 = (n_580 ^ (csa_tree_add_106_2_groupi_n_818 ^ n_190));
 assign csa_tree_add_106_2_groupi_n_886 = ~(n_542 ^ n_56);
 assign csa_tree_add_106_2_groupi_n_0 = ~((n_540 & (n_541 & n_411)) | (n_547 & n_1477));
 assign n_556 = ~((n_577 & n_465) | (n_557 & stall));
 assign n_545 = ((n_839 & n_597) | ((n_597 & n_64) | (n_64 & n_839)));
 assign csa_tree_add_106_2_groupi_n_693 = (n_597 ^ (n_64 ^ n_839));
 assign n_555 = ((n_316 & n_603) | ((n_603 & n_799) | (n_799 & n_316)));
 assign n_554 = (n_603 ^ (n_799 ^ n_316));
 assign csa_tree_add_106_2_groupi_n_870 = ((n_813 & n_618) | ((n_618 & n_80) | (n_80 & n_813)));
 assign n_551 = (n_618 ^ (n_80 ^ n_813));
 assign csa_tree_add_106_2_groupi_n_1087 = ((n_1003 & n_608) | ((n_608 & n_557) | (n_557 & n_1003)));
 assign csa_tree_add_106_2_groupi_n_1088 = (n_608 ^ (n_557 ^ n_1003));
 assign csa_tree_add_106_2_groupi_n_982 = ((n_38 & n_172) | ((n_172 & n_58) | (n_58 & n_38)));
 assign n_550 = (n_172 ^ (n_58 ^ n_38));
 assign csa_tree_add_106_2_groupi_n_880 = ((n_836 & n_599) | ((n_599 & n_85) | (n_85 & n_836)));
 assign csa_tree_add_106_2_groupi_n_881 = (n_599 ^ (n_85 ^ n_836));
 assign csa_tree_add_106_2_groupi_n_995 = ((n_59 & n_609) | ((n_609 & n_39) | (n_39 & n_59)));
 assign csa_tree_add_106_2_groupi_n_996 = (n_609 ^ (n_39 ^ n_59));
 assign csa_tree_add_92_2_groupi_n_188 = ((n_338 & n_1366) | ((n_1366 & n_335) | (n_335 & n_338)));
 assign csa_tree_add_92_2_groupi_n_189 = (n_1366 ^ (n_335 ^ n_338));
 assign csa_tree_add_106_2_groupi_n_958 = ((n_814 & n_611) | ((n_611 & n_353) | (n_353 & n_814)));
 assign csa_tree_add_106_2_groupi_n_959 = (n_611 ^ (n_353 ^ n_814));
 assign csa_tree_add_106_2_groupi_n_364 = ~((n_571 | n_412) & (n_680 | n_414));
 assign csa_tree_add_106_2_groupi_n_446 = ~((n_569 | n_378) & (n_677 | n_380));
 assign csa_tree_add_106_2_groupi_n_451 = ~((n_569 | n_380) & (n_1083 | n_378));
 assign csa_tree_add_106_2_groupi_n_521 = ~((n_572 | n_391) & (n_1097 | n_389));
 assign csa_tree_add_106_2_groupi_n_583 = ~((n_570 | n_399) & (n_1101 | n_397));
 assign csa_tree_add_106_2_groupi_n_515 = ~((n_572 | n_389) & (n_678 | n_391));
 assign csa_tree_add_106_2_groupi_n_578 = ~((n_570 | n_397) & (n_679 | n_399));
 assign csa_tree_add_106_2_groupi_n_369 = ~((n_571 | n_414) & (n_1114 | n_412));
 assign csa_tree_add_86_2_n_954 = ((n_789 & n_718) | ((n_718 & n_125) | (n_125 & n_789)));
 assign csa_tree_add_86_2_n_955 = (n_718 ^ (n_125 ^ n_789));
 assign n_577 = ((n_667 & csa_tree_add_106_2_groupi_n_976) | ((csa_tree_add_106_2_groupi_n_976 & csa_tree_add_106_2_groupi_n_888)
    | (csa_tree_add_106_2_groupi_n_888 & n_667)));
 assign n_576 = (csa_tree_add_106_2_groupi_n_976 ^ (csa_tree_add_106_2_groupi_n_888 ^ n_667));
 assign n_564 = ((csa_tree_add_92_2_groupi_n_182 & n_590) | ((n_590 & n_989) | (n_989 & csa_tree_add_92_2_groupi_n_182)));
 assign n_563 = (n_590 ^ (n_989 ^ csa_tree_add_92_2_groupi_n_182));
 assign n_596 = ((n_703 & csa_tree_add_106_2_groupi_n_370) | ((csa_tree_add_106_2_groupi_n_370 & csa_tree_add_106_2_groupi_n_718)
    | (csa_tree_add_106_2_groupi_n_718 & n_703)));
 assign n_595 = (csa_tree_add_106_2_groupi_n_370 ^ (csa_tree_add_106_2_groupi_n_718 ^ n_703));
 assign n_566 = ((n_328 & n_178) | ((n_178 & n_1400) | (n_1400 & n_328)));
 assign n_565 = (n_178 ^ (n_1400 ^ n_328));
 assign n_591 = ~n_601;
 assign n_594 = ~(n_176 | ~(n_438 | n_465));
 assign n_573 = ((n_62 & ~n_465) | (n_592 & n_465));
 assign n_601 = ~((csa_tree_mul_77_11_groupi_n_408 | (n_177 | stall)) & (n_343 | n_465));
 assign mul_109_11_n_630 = ~(mul_109_11_n_28 | ((n_1457 & n_1458) | (mul_109_11_n_2 & n_362)));
 assign n_542 = ~((n_574 | n_379) & (n_600 | n_381));
 assign n_543 = ~((n_544 | n_413) & (n_598 | n_415));
 assign n_534 = ~((n_544 | n_415) & (n_546 | n_413));
 assign n_659 = ((n_959 & n_1014) | ((n_1014 & n_108) | (n_108 & n_959)));
 assign n_658 = (n_1014 ^ (n_108 ^ n_959));
 assign n_579 = ((n_187 & n_1041) | ((n_1041 & csa_tree_add_106_2_groupi_n_872) | (csa_tree_add_106_2_groupi_n_872
    & n_187)));
 assign n_578 = (n_1041 ^ (csa_tree_add_106_2_groupi_n_872 ^ n_187));
 assign n_581 = ((n_237 & n_1045) | ((n_1045 & n_695) | (n_695 & n_237)));
 assign n_580 = (n_1045 ^ (n_695 ^ n_237));
 assign csa_tree_add_106_2_groupi_n_968 = ((n_844 & n_607) | ((n_607 & n_314) | (n_314 & n_844)));
 assign csa_tree_add_106_2_groupi_n_969 = (n_607 ^ (n_314 ^ n_844));
 assign csa_tree_add_92_2_groupi_n_194 = ((n_336 & n_1398) | ((n_1398 & n_333) | (n_333 & n_336)));
 assign csa_tree_add_92_2_groupi_n_195 = (n_1398 ^ (n_333 ^ n_336));
 assign n_176 = ~(stall | (csa_tree_mul_77_11_groupi_n_408 & n_177));
 assign n_593 = ~((n_180 & n_465) | (n_797 & stall));
 assign n_540 = ~(n_548 & n_417);
 assign n_541 = ~(n_549 & n_419);
 assign n_570 = ~((n_1426 & n_402) | (csa_tree_add_106_2_groupi_n_49 & n_160));
 assign n_572 = ~((n_1426 & n_395) | (csa_tree_add_106_2_groupi_n_49 & n_393));
 assign n_569 = ~((n_1426 & n_384) | (csa_tree_add_106_2_groupi_n_49 & n_382));
 assign n_571 = ~((n_1426 & n_418) | (csa_tree_add_106_2_groupi_n_49 & n_416));
 assign n_568 = ((n_1375 & csa_tree_add_92_2_groupi_n_149) | ((csa_tree_add_92_2_groupi_n_149 & n_196)
    | (n_196 & n_1375)));
 assign n_567 = (csa_tree_add_92_2_groupi_n_149 ^ (n_196 ^ n_1375));
 assign n_661 = ((n_1374 & n_1404) | ((n_1404 & n_936) | (n_936 & n_1374)));
 assign n_660 = (n_1404 ^ (n_936 ^ n_1374));
 assign csa_tree_add_86_2_n_940 = ((n_262 & n_788) | ((n_788 & n_157) | (n_157 & n_262)));
 assign csa_tree_add_86_2_n_941 = (n_788 ^ (n_157 ^ n_262));
 assign n_583 = ((csa_tree_add_86_2_n_436 & csa_tree_add_86_2_n_920) | ((csa_tree_add_86_2_n_920 & n_700)
    | (n_700 & csa_tree_add_86_2_n_436)));
 assign n_582 = (csa_tree_add_86_2_n_920 ^ (n_700 ^ csa_tree_add_86_2_n_436));
 assign n_663 = ((n_979 & csa_tree_add_106_2_groupi_n_558) | ((csa_tree_add_106_2_groupi_n_558 & n_951)
    | (n_951 & n_979)));
 assign n_662 = (csa_tree_add_106_2_groupi_n_558 ^ (n_951 ^ n_979));
 assign n_546 = ~n_547;
 assign n_548 = ~n_549;
 assign csa_tree_mul_77_11_groupi_n_619 = (n_584 & n_340);
 assign n_574 = ~((n_383 & ~n_575) | (n_385 & n_575));
 assign n_592 = ~(n_681 ^ csa_tree_add_106_2_groupi_n_855);
 assign csa_tree_add_106_2_groupi_n_821 = ~(n_617 ^ n_102);
 assign n_544 = ~((n_417 & ~n_575) | (n_419 & n_575));
 assign n_547 = ~(n_588 ^ n_417);
 assign csa_tree_add_106_2_groupi_n_3 = ~(csa_tree_add_106_2_groupi_n_222 & ~csa_tree_add_106_2_groupi_n_218);
 assign n_549 = ~(n_587 ^ n_7);
 assign final_adder_add_86_2_n_19 = ((n_1148 & n_657) | ((n_657 & n_442) | (n_442 & n_1148)));
 assign n_1426 = (n_657 ^ (n_442 ^ n_1148));
 assign n_664 = ((n_32 & n_1009) | ((n_1009 & n_28) | (n_28 & n_32)));
 assign n_1457 = (n_1009 ^ (n_28 ^ n_32));
 assign n_707 = ((n_929 & csa_tree_add_86_2_n_921) | ((csa_tree_add_86_2_n_921 & csa_tree_add_86_2_n_903)
    | (csa_tree_add_86_2_n_903 & n_929)));
 assign n_706 = (csa_tree_add_86_2_n_921 ^ (csa_tree_add_86_2_n_903 ^ n_929));
 assign n_668 = ((n_1019 & n_1032) | ((n_1032 & csa_tree_add_106_2_groupi_n_810) | (csa_tree_add_106_2_groupi_n_810
    & n_1019)));
 assign n_667 = (n_1032 ^ (csa_tree_add_106_2_groupi_n_810 ^ n_1019));
 assign n_612 = ((n_807 & n_833) | ((n_833 & n_315) | (n_315 & n_807)));
 assign csa_tree_add_106_2_groupi_n_931 = (n_833 ^ (n_315 ^ n_807));
 assign n_670 = ((csa_tree_add_86_2_n_891 & csa_tree_add_86_2_n_871) | ((csa_tree_add_86_2_n_871 & n_988)
    | (n_988 & csa_tree_add_86_2_n_891)));
 assign n_669 = (csa_tree_add_86_2_n_871 ^ (n_988 ^ csa_tree_add_86_2_n_891));
 assign n_672 = ((n_239 & n_1023) | ((n_1023 & n_1011) | (n_1011 & n_239)));
 assign n_671 = (n_1023 ^ (n_1011 ^ n_239));
 assign csa_tree_add_92_2_groupi_n_208 = ((n_332 & n_1369) | ((n_1369 & n_330) | (n_330 & n_332)));
 assign n_178 = (n_1369 ^ (n_330 ^ n_332));
 assign csa_tree_add_92_2_groupi_n_198 = ((n_334 & n_1368) | ((n_1368 & n_331) | (n_331 & n_334)));
 assign csa_tree_add_92_2_groupi_n_199 = (n_1368 ^ (n_331 ^ n_334));
 assign n_177 = ((n_996 & csa_tree_mul_77_11_groupi_n_335) | ((csa_tree_mul_77_11_groupi_n_335 & csa_tree_mul_77_11_groupi_n_330)
    | (csa_tree_mul_77_11_groupi_n_330 & n_996)));
 assign n_693 = (csa_tree_mul_77_11_groupi_n_335 ^ (csa_tree_mul_77_11_groupi_n_330 ^ n_996));
 assign n_180 = ((csa_tree_mul_77_11_groupi_n_298 & n_957) | ((n_957 & csa_tree_mul_77_11_groupi_n_249)
    | (csa_tree_mul_77_11_groupi_n_249 & csa_tree_mul_77_11_groupi_n_298)));
 assign n_179 = (n_957 ^ (csa_tree_mul_77_11_groupi_n_249 ^ csa_tree_mul_77_11_groupi_n_298));
 assign n_584 = ~(n_339 & (n_175 | csa_tree_mul_77_11_groupi_n_514));
 assign n_682 = ~((csa_tree_add_106_2_groupi_n_336 & n_465) | (n_1178 & stall));
 assign n_708 = ~((n_782 & (n_1353 & n_465)) | (n_709 & stall));
 assign n_613 = ~((n_675 | csa_tree_add_106_2_groupi_n_230) & (csa_tree_add_106_2_groupi_n_61 | csa_tree_add_106_2_groupi_n_336));
 assign n_673 = (n_684 ^ n_674);
 assign n_614 = ~((csa_tree_add_106_2_groupi_n_230 & n_465) | (n_1179 & stall));
 assign mul_109_11_n_520 = ~((n_586 | n_311) & (n_719 | n_585));
 assign n_615 = ~((n_705 & n_465) | (n_791 & stall));
 assign n_616 = ~((n_704 & n_465) | (n_250 & stall));
 assign mul_109_11_n_521 = ~((n_586 | n_585) & (n_750 | n_311));
 assign csa_tree_add_106_2_groupi_n_262 = ~((n_710 | n_1437) & (n_675 | csa_tree_add_106_2_groupi_n_38));
 assign csa_tree_add_106_2_groupi_n_222 = ~(csa_tree_add_106_2_groupi_n_36 ^ csa_tree_add_106_2_groupi_n_38);
 assign csa_tree_add_86_2_n_956 = ((n_139 & n_787) | ((n_787 & n_127) | (n_127 & n_139)));
 assign csa_tree_add_86_2_n_957 = (n_787 ^ (n_127 ^ n_139));
 assign csa_tree_add_106_2_groupi_n_675 = ((n_236 & n_846) | ((n_846 & n_132) | (n_132 & n_236)));
 assign csa_tree_add_106_2_groupi_n_676 = (n_846 ^ (n_132 ^ n_236));
 assign n_603 = ((n_368 & n_808) | ((n_808 & n_169) | (n_169 & n_368)));
 assign n_602 = (n_808 ^ (n_169 ^ n_368));
 assign n_605 = ((n_386 & n_810) | ((n_810 & n_134) | (n_134 & n_386)));
 assign n_604 = (n_810 ^ (n_134 ^ n_386));
 assign csa_tree_add_106_2_groupi_n_954 = ((n_42 & n_827) | ((n_827 & n_35) | (n_35 & n_42)));
 assign csa_tree_add_106_2_groupi_n_955 = (n_827 ^ (n_35 ^ n_42));
 assign n_182 = ((csa_tree_add_106_2_groupi_n_805 & n_1027) | ((n_1027 & n_238) | (n_238 & csa_tree_add_106_2_groupi_n_805)));
 assign n_181 = (n_1027 ^ (n_238 ^ csa_tree_add_106_2_groupi_n_805));
 assign n_184 = ((n_1043 & n_1018) | ((n_1018 & csa_tree_add_106_2_groupi_n_806) | (csa_tree_add_106_2_groupi_n_806
    & n_1043)));
 assign n_183 = (n_1018 ^ (csa_tree_add_106_2_groupi_n_806 ^ n_1043));
 assign n_186 = ((csa_tree_add_106_2_groupi_n_809 & n_1026) | ((n_1026 & csa_tree_add_106_2_groupi_n_738)
    | (csa_tree_add_106_2_groupi_n_738 & csa_tree_add_106_2_groupi_n_809)));
 assign n_185 = (n_1026 ^ (csa_tree_add_106_2_groupi_n_738 ^ csa_tree_add_106_2_groupi_n_809));
 assign n_188 = ((csa_tree_add_106_2_groupi_n_807 & n_1030) | ((n_1030 & csa_tree_add_106_2_groupi_n_742)
    | (csa_tree_add_106_2_groupi_n_742 & csa_tree_add_106_2_groupi_n_807)));
 assign n_187 = (n_1030 ^ (csa_tree_add_106_2_groupi_n_742 ^ csa_tree_add_106_2_groupi_n_807));
 assign csa_tree_add_106_2_groupi_n_797 = ((n_1065 & n_847) | ((n_847 & n_161) | (n_161 & n_1065)));
 assign csa_tree_add_106_2_groupi_n_798 = (n_847 ^ (n_161 ^ n_1065));
 assign n_190 = ((csa_tree_add_106_2_groupi_n_824 & n_1022) | ((n_1022 & csa_tree_add_106_2_groupi_n_750)
    | (csa_tree_add_106_2_groupi_n_750 & csa_tree_add_106_2_groupi_n_824)));
 assign n_189 = (n_1022 ^ (csa_tree_add_106_2_groupi_n_750 ^ csa_tree_add_106_2_groupi_n_824));
 assign n_192 = ((n_240 & n_1020) | ((n_1020 & csa_tree_add_106_2_groupi_n_817) | (csa_tree_add_106_2_groupi_n_817
    & n_240)));
 assign n_191 = (n_1020 ^ (csa_tree_add_106_2_groupi_n_817 ^ n_240));
 assign n_194 = ((n_1062 & n_1058) | ((n_1058 & csa_tree_add_106_2_groupi_n_825) | (csa_tree_add_106_2_groupi_n_825
    & n_1062)));
 assign n_193 = (n_1058 ^ (csa_tree_add_106_2_groupi_n_825 ^ n_1062));
 assign csa_tree_add_106_2_groupi_n_852 = ((n_352 & n_826) | ((n_826 & n_103) | (n_103 & n_352)));
 assign csa_tree_add_106_2_groupi_n_853 = (n_826 ^ (n_103 ^ n_352));
 assign csa_tree_add_106_2_groupi_n_932 = ((n_805 & n_842) | ((n_842 & n_313) | (n_313 & n_805)));
 assign csa_tree_add_106_2_groupi_n_933 = (n_842 ^ (n_313 ^ n_805));
 assign n_607 = ((n_816 & n_812) | ((n_812 & n_168) | (n_168 & n_816)));
 assign n_606 = (n_812 ^ (n_168 ^ n_816));
 assign n_609 = ((n_46 & n_829) | ((n_829 & n_41) | (n_41 & n_46)));
 assign n_608 = (n_829 ^ (n_41 ^ n_46));
 assign n_611 = ((n_323 & n_848) | ((n_848 & n_162) | (n_162 & n_323)));
 assign csa_tree_add_106_2_groupi_n_921 = (n_848 ^ (n_162 ^ n_323));
 assign csa_tree_add_106_2_groupi_n_936 = ((n_63 & n_806) | ((n_806 & n_47) | (n_47 & n_63)));
 assign n_610 = (n_806 ^ (n_47 ^ n_63));
 assign n_1366 = ((n_126 & n_942) | ((n_942 & n_123) | (n_123 & n_126)));
 assign n_1398 = (n_942 ^ (n_123 ^ n_126));
 assign n_587 = ~((n_589 & n_1462) | (n_4 & n_3));
 assign n_681 = ~((n_783 | n_398) & (n_1025 | n_399));
 assign n_575 = ~(n_676 ^ n_5);
 assign csa_tree_add_106_2_groupi_n_436 = ~((n_677 | n_378) & (n_886 | n_380));
 assign csa_tree_add_106_2_groupi_n_499 = ~((n_678 | n_389) & (n_891 | n_391));
 assign csa_tree_add_106_2_groupi_n_573 = ~((n_679 | n_397) & (n_896 | n_399));
 assign csa_tree_add_106_2_groupi_n_367 = ~((n_680 | n_412) & (n_900 | n_414));
 assign n_588 = ~(n_589 ^ csa_tree_add_92_2_groupi_n_65);
 assign n_617 = ~((n_711 | n_390) & (n_837 | n_392));
 assign n_597 = ~((n_598 | n_413) & (n_173 | n_415));
 assign n_618 = ~((n_619 | n_379) & (n_840 | n_381));
 assign n_172 = ~((n_173 | n_413) & (n_828 | n_415));
 assign n_599 = ~((n_600 | n_379) & (n_619 | n_381));
 assign csa_tree_add_106_2_groupi_n_38 = ~n_1437;
 assign n_196 = ((csa_tree_add_92_2_groupi_n_99 & n_1376) | ((n_1376 & n_944) | (n_944 & csa_tree_add_92_2_groupi_n_99)));
 assign n_195 = (n_1376 ^ (n_944 ^ csa_tree_add_92_2_groupi_n_99));
 assign n_699 = ((n_985 & csa_tree_add_106_2_groupi_n_977) | ((csa_tree_add_106_2_groupi_n_977 & csa_tree_add_106_2_groupi_n_1018)
    | (csa_tree_add_106_2_groupi_n_1018 & n_985)));
 assign n_698 = (csa_tree_add_106_2_groupi_n_977 ^ (csa_tree_add_106_2_groupi_n_1018 ^ n_985));
 assign n_701 = ((n_954 & csa_tree_add_86_2_n_125) | ((csa_tree_add_86_2_n_125 & csa_tree_add_86_2_n_192)
    | (csa_tree_add_86_2_n_192 & n_954)));
 assign n_700 = (csa_tree_add_86_2_n_125 ^ (csa_tree_add_86_2_n_192 ^ n_954));
 assign n_198 = ((csa_tree_add_86_2_n_902 & csa_tree_add_86_2_n_158) | ((csa_tree_add_86_2_n_158 & n_967)
    | (n_967 & csa_tree_add_86_2_n_902)));
 assign n_197 = (csa_tree_add_86_2_n_158 ^ (n_967 ^ csa_tree_add_86_2_n_902));
 assign n_697 = ((n_993 & csa_tree_add_86_2_n_105) | ((csa_tree_add_86_2_n_105 & csa_tree_add_86_2_n_154)
    | (csa_tree_add_86_2_n_154 & n_993)));
 assign n_696 = (csa_tree_add_86_2_n_105 ^ (csa_tree_add_86_2_n_154 ^ n_993));
 assign n_200 = ((csa_tree_add_106_2_groupi_n_504 & n_937) | ((n_937 & csa_tree_add_106_2_groupi_n_770)
    | (csa_tree_add_106_2_groupi_n_770 & csa_tree_add_106_2_groupi_n_504)));
 assign n_199 = (n_937 ^ (csa_tree_add_106_2_groupi_n_770 ^ csa_tree_add_106_2_groupi_n_504));
 assign n_666 = ((csa_tree_add_106_2_groupi_n_465 & csa_tree_add_106_2_groupi_n_779) | ((csa_tree_add_106_2_groupi_n_779
    & n_933) | (n_933 & csa_tree_add_106_2_groupi_n_465)));
 assign n_665 = (csa_tree_add_106_2_groupi_n_779 ^ (n_933 ^ csa_tree_add_106_2_groupi_n_465));
 assign n_705 = ((n_934 & csa_tree_mul_77_11_groupi_n_346) | ((csa_tree_mul_77_11_groupi_n_346 & csa_tree_mul_77_11_groupi_n_401)
    | (csa_tree_mul_77_11_groupi_n_401 & n_934)));
 assign n_704 = (csa_tree_mul_77_11_groupi_n_346 ^ (csa_tree_mul_77_11_groupi_n_401 ^ n_934));
 assign n_590 = ((csa_tree_add_86_2_n_887 & n_926) | ((n_926 & csa_tree_add_86_2_n_894) | (csa_tree_add_86_2_n_894
    & csa_tree_add_86_2_n_887)));
 assign n_654 = (n_926 ^ (csa_tree_add_86_2_n_894 ^ csa_tree_add_86_2_n_887));
 assign n_703 = ((csa_tree_add_106_2_groupi_n_661 & csa_tree_add_106_2_groupi_n_362) | ((csa_tree_add_106_2_groupi_n_362
    & n_1172) | (n_1172 & csa_tree_add_106_2_groupi_n_661)));
 assign n_702 = (csa_tree_add_106_2_groupi_n_362 ^ (n_1172 ^ csa_tree_add_106_2_groupi_n_661));
 assign final_adder_add_69_2_n_2 = (({in2[1]} & n_274) | ((n_274 & {in1[1]}) | ({in1[1]} & {in2[1]})));
 assign n_1437 = (n_274 ^ ({in1[1]} ^ {in2[1]}));
 assign n_656 = ((n_110 & n_329) | ((n_329 & n_657) | (n_657 & n_110)));
 assign n_655 = (n_329 ^ (n_657 ^ n_110));
 assign n_685 = ~n_714;
 assign n_714 = ~((csa_tree_mul_77_11_groupi_n_452 | (n_794 | stall)) & (n_150 | n_465));
 assign mul_109_11_n_365 = ~(n_174 ^ n_310);
 assign mul_109_11_n_246 = ~(n_174 ^ n_88);
 assign n_683 = ~(n_781 & ~(n_684 & n_1353));
 assign n_175 = (csa_tree_mul_77_11_groupi_n_487 & (csa_tree_mul_77_11_groupi_n_590 | csa_tree_mul_77_11_groupi_n_606));
 assign n_688 = ~(n_690 & (n_689 | n_223));
 assign csa_tree_add_106_2_groupi_n_233 = ~((n_710 | n_1435) & (n_675 | csa_tree_add_106_2_groupi_n_39));
 assign n_586 = ~(n_174 ^ n_136);
 assign csa_tree_mul_77_11_groupi_n_514 = (n_691 | n_438);
 assign csa_tree_add_106_2_groupi_n_177 = ~((n_710 | n_1433) & (n_675 | csa_tree_add_106_2_groupi_n_7));
 assign csa_tree_add_106_2_groupi_n_2 = ~(csa_tree_add_106_2_groupi_n_223 & ~csa_tree_add_106_2_groupi_n_215);
 assign csa_tree_add_106_2_groupi_n_4 = ~(csa_tree_add_106_2_groupi_n_221 & ~csa_tree_add_106_2_groupi_n_217);
 assign csa_tree_add_106_2_groupi_n_344 = ~(csa_tree_add_106_2_groupi_n_225 & ~csa_tree_add_106_2_groupi_n_211);
 assign csa_tree_add_86_2_n_912 = ((n_273 & n_275) | ((n_275 & n_141) | (n_141 & n_273)));
 assign n_789 = (n_275 ^ (n_141 ^ n_273));
 assign csa_tree_add_86_2_n_906 = ((n_267 & n_276) | ((n_276 & n_142) | (n_142 & n_267)));
 assign csa_tree_add_86_2_n_907 = (n_276 ^ (n_142 ^ n_267));
 assign csa_tree_add_86_2_n_896 = ((n_268 & n_272) | ((n_272 & n_155) | (n_155 & n_268)));
 assign csa_tree_add_86_2_n_897 = (n_272 ^ (n_155 ^ n_268));
 assign csa_tree_add_86_2_n_918 = ((n_156 & n_271) | ((n_271 & n_261) | (n_261 & n_156)));
 assign csa_tree_add_86_2_n_919 = (n_271 ^ (n_261 ^ n_156));
 assign csa_tree_add_86_2_n_876 = ((n_1383 & n_158) | ((n_158 & n_1430) | (n_1430 & n_1383)));
 assign csa_tree_add_86_2_n_877 = (n_158 ^ (n_1430 ^ n_1383));
 assign csa_tree_add_86_2_n_872 = ((n_270 & n_159) | ((n_159 & n_260) | (n_260 & n_270)));
 assign csa_tree_add_86_2_n_873 = (n_159 ^ (n_260 ^ n_270));
 assign n_695 = ((csa_tree_add_106_2_groupi_n_689 & n_241) | ((n_241 & csa_tree_add_106_2_groupi_n_776)
    | (csa_tree_add_106_2_groupi_n_776 & csa_tree_add_106_2_groupi_n_689)));
 assign n_694 = (n_241 ^ (csa_tree_add_106_2_groupi_n_776 ^ csa_tree_add_106_2_groupi_n_689));
 assign csa_tree_add_86_2_n_608 = ((n_266 & n_1378) | ((n_1378 & n_115) | (n_115 & n_266)));
 assign csa_tree_add_86_2_n_609 = (n_1378 ^ (n_115 ^ n_266));
 assign csa_tree_mul_77_11_groupi_n_503 = ~(n_792 & n_791);
 assign n_778 = ~(n_1379 ^ n_1351);
 assign n_779 = ~(n_780 ^ n_222);
 assign n_781 = ~(n_782 & (n_684 | n_1353));
 assign n_691 = ~(csa_tree_mul_77_11_groupi_n_460 | ~n_343);
 assign csa_tree_mul_77_11_groupi_n_499 = ~(n_792 | n_791);
 assign n_679 = ~((n_1427 & n_402) | (csa_tree_add_106_2_groupi_n_53 & n_160));
 assign n_680 = ~((n_1427 & n_418) | (csa_tree_add_106_2_groupi_n_53 & n_416));
 assign csa_tree_mul_77_11_groupi_n_487 = ~(csa_tree_mul_77_11_groupi_n_459 | ~n_343);
 assign n_173 = ~((n_419 & ~n_716) | (n_417 & n_716));
 assign n_598 = ~((n_419 & ~n_692) | (n_417 & n_692));
 assign csa_tree_add_106_2_groupi_n_248 = ~((n_1446 & ~n_1346) | (csa_tree_add_106_2_groupi_n_40 & n_1346));
 assign n_677 = ~((n_1427 & n_384) | (csa_tree_add_106_2_groupi_n_53 & n_382));
 assign n_678 = ~((n_1427 & n_395) | (csa_tree_add_106_2_groupi_n_53 & n_393));
 assign n_619 = ~((n_385 & ~n_716) | (n_383 & n_716));
 assign n_589 = ~(n_686 & ~csa_tree_add_92_2_groupi_n_89);
 assign csa_tree_add_106_2_groupi_n_230 = ~(csa_tree_add_106_2_groupi_n_336 & (n_1431 | n_796));
 assign mul_109_11_n_114 = ~((n_1458 | n_96) & (mul_109_11_n_43 | n_746));
 assign n_711 = ~((n_396 & ~n_716) | (n_394 & n_716));
 assign n_713 = ~((csa_tree_add_106_2_groupi_n_228 & n_465) | (n_203 & stall));
 assign n_785 = ~((n_962 & n_465) | (n_251 & stall));
 assign n_784 = ~((n_995 & n_465) | (n_798 & stall));
 assign n_790 = ~((csa_tree_add_106_2_groupi_n_338 & n_465) | (n_202 & stall));
 assign mul_109_11_n_82 = ~((n_1458 | n_362) & (mul_109_11_n_43 | mul_109_11_n_38));
 assign mul_109_11_n_88 = ~((n_106 | n_1458) & (mul_109_11_n_43 | n_749));
 assign mul_109_11_n_89 = ~((n_1458 | n_1) & (mul_109_11_n_43 | n_751));
 assign mul_109_11_n_90 = ~((n_1458 | n_433) & (mul_109_11_n_43 | n_777));
 assign mul_109_11_n_99 = ~((n_1458 | n_90) & (mul_109_11_n_43 | n_743));
 assign mul_109_11_n_98 = ~((n_1458 | n_92) & (mul_109_11_n_43 | n_744));
 assign mul_109_11_n_113 = ~((n_1458 | n_95) & (mul_109_11_n_43 | n_745));
 assign mul_109_11_n_238 = ~((mul_109_11_n_43 & ~n_45) | (n_1458 & n_45));
 assign mul_109_11_n_125 = ~((n_1458 | n_97) & (mul_109_11_n_43 | n_747));
 assign mul_109_11_n_124 = ~((n_1458 | n_98) & (mul_109_11_n_43 | n_748));
 assign n_783 = ((n_402 & ~n_717) | (n_160 & n_717));
 assign mul_109_11_n_148 = ~((n_1458 | n_99) & (mul_109_11_n_43 | n_1198));
 assign mul_109_11_n_78 = ~((n_1458 | n_100) & (mul_109_11_n_43 | n_1197));
 assign n_600 = ~((n_385 & ~n_692) | (n_383 & n_692));
 assign csa_tree_add_106_2_groupi_n_113 = ~((n_1428 | n_1431) & (csa_tree_add_106_2_groupi_n_61 | csa_tree_add_106_2_groupi_n_44));
 assign n_676 = ~(n_687 ^ n_9);
 assign csa_tree_add_106_2_groupi_n_221 = ~(csa_tree_add_106_2_groupi_n_73 ^ csa_tree_add_106_2_groupi_n_40);
 assign csa_tree_add_106_2_groupi_n_223 = ~(csa_tree_add_106_2_groupi_n_74 ^ csa_tree_add_106_2_groupi_n_39);
 assign csa_tree_add_106_2_groupi_n_225 = ~(csa_tree_add_106_2_groupi_n_37 ^ csa_tree_add_106_2_groupi_n_7);
 assign n_674 = (n_782 ^ n_1353);
 assign n_675 = ~n_710;
 assign n_959 = ((n_107 & n_109) | ((n_109 & n_93) | (n_93 & n_107)));
 assign n_958 = (n_109 ^ (n_93 ^ n_107));
 assign csa_tree_add_86_2_n_964 = ((n_128 & n_146) | ((n_146 & n_140) | (n_140 & n_128)));
 assign n_942 = (n_146 ^ (n_140 ^ n_128));
 assign csa_tree_add_106_2_groupi_n_989 = ((n_36 & n_43) | ((n_43 & n_21) | (n_21 & n_36)));
 assign n_1003 = (n_43 ^ (n_21 ^ n_36));
 assign n_936 = ((n_1405 & n_1375) | ((n_1375 & final_adder_add_86_2_n_3) | (final_adder_add_86_2_n_3
    & n_1405)));
 assign n_710 = (n_1375 ^ (final_adder_add_86_2_n_3 ^ n_1405));
 assign n_788 = ((n_356 & n_269) | ((n_269 & n_143) | (n_143 & n_356)));
 assign n_787 = (n_269 ^ (n_143 ^ n_356));
 assign csa_tree_add_92_2_groupi_n_276 = ((n_30 & n_709) | ((n_709 & n_852) | (n_852 & n_30)));
 assign n_174 = (n_709 ^ (n_852 ^ n_30));
 assign csa_tree_mul_77_11_groupi_n_469 = ((n_167 & n_346) | ((n_346 & n_165) | (n_165 & n_167)));
 assign n_792 = (n_346 ^ (n_165 ^ n_167));
 assign csa_tree_add_86_2_n_668 = ((n_116 & n_263) | ((n_263 & n_354) | (n_354 & n_116)));
 assign n_718 = (n_263 ^ (n_354 ^ n_116));
 assign csa_tree_add_106_2_groupi_n_1073 = ((n_22 & n_25) | ((n_25 & n_16) | (n_16 & n_22)));
 assign n_974 = (n_25 ^ (n_16 ^ n_22));
 assign n_1367 = ((n_144 & n_147) | ((n_147 & n_124) | (n_124 & n_144)));
 assign n_1399 = (n_147 ^ (n_124 ^ n_144));
 assign n_793 = ~(csa_tree_mul_77_11_groupi_n_452 & n_794);
 assign csa_tree_mul_77_11_groupi_n_460 = ~(n_786 & n_373);
 assign n_690 = ~(n_780 & n_1370);
 assign n_689 = ~(n_780 | n_1370);
 assign csa_tree_add_106_2_groupi_n_336 = ~(n_1431 & n_796);
 assign csa_tree_add_106_2_groupi_n_539 = ~(n_437 & (n_715 | n_429));
 assign n_795 = ~(n_1446 & n_1447);
 assign mul_109_11_n_547 = ~((n_1151 & (n_1165 & n_370)) | (mul_109_11_n_348 & mul_109_11_n_383));
 assign n_686 = ~(n_687 & (n_5 | n_9));
 assign csa_tree_add_106_2_groupi_n_586 = ~((n_715 | n_78) & (n_821 | n_429));
 assign csa_tree_add_106_2_groupi_n_628 = ~((n_712 | n_424) & (n_423 | n_439));
 assign csa_tree_add_106_2_groupi_n_598 = ~((n_712 | n_423) & (n_1494 | n_424));
 assign csa_tree_mul_77_11_groupi_n_459 = ~(n_786 | n_373);
 assign csa_tree_add_106_2_groupi_n_39 = ~n_1435;
 assign csa_tree_add_106_2_groupi_n_44 = ~n_1431;
 assign csa_tree_add_106_2_groupi_n_40 = ~n_1446;
 assign csa_tree_add_106_2_groupi_n_7 = ~n_1433;
 assign n_986 = ((csa_tree_add_106_2_groupi_n_889 & csa_tree_add_106_2_groupi_n_974) | ((csa_tree_add_106_2_groupi_n_974
    & csa_tree_add_106_2_groupi_n_924) | (csa_tree_add_106_2_groupi_n_924 & csa_tree_add_106_2_groupi_n_889)));
 assign n_985 = (csa_tree_add_106_2_groupi_n_974 ^ (csa_tree_add_106_2_groupi_n_924 ^ csa_tree_add_106_2_groupi_n_889));
 assign n_946 = ((csa_tree_add_86_2_n_870 & csa_tree_add_86_2_n_437) | ((csa_tree_add_86_2_n_437 & csa_tree_add_86_2_n_890)
    | (csa_tree_add_86_2_n_890 & csa_tree_add_86_2_n_870)));
 assign n_945 = (csa_tree_add_86_2_n_437 ^ (csa_tree_add_86_2_n_890 ^ csa_tree_add_86_2_n_870));
 assign csa_tree_add_92_2_groupi_n_164 = ((n_408 & n_1365) | ((n_1365 & n_337) | (n_337 & n_408)));
 assign csa_tree_add_92_2_groupi_n_165 = (n_1365 ^ (n_337 ^ n_408));
 assign n_1007 = ((csa_tree_add_106_2_groupi_n_1019 & csa_tree_add_106_2_groupi_n_975) | ((csa_tree_add_106_2_groupi_n_975
    & csa_tree_add_106_2_groupi_n_1005) | (csa_tree_add_106_2_groupi_n_1005 & csa_tree_add_106_2_groupi_n_1019)));
 assign n_1006 = (csa_tree_add_106_2_groupi_n_975 ^ (csa_tree_add_106_2_groupi_n_1005 ^ csa_tree_add_106_2_groupi_n_1019));
 assign n_951 = ((csa_tree_add_106_2_groupi_n_631 & csa_tree_add_106_2_groupi_n_563) | ((csa_tree_add_106_2_groupi_n_563
    & csa_tree_add_106_2_groupi_n_686) | (csa_tree_add_106_2_groupi_n_686 & csa_tree_add_106_2_groupi_n_631)));
 assign n_950 = (csa_tree_add_106_2_groupi_n_563 ^ (csa_tree_add_106_2_groupi_n_686 ^ csa_tree_add_106_2_groupi_n_631));
 assign n_931 = ((csa_tree_mul_77_11_groupi_n_324 & csa_tree_mul_77_11_groupi_n_345) | ((csa_tree_mul_77_11_groupi_n_345
    & csa_tree_mul_77_11_groupi_n_299) | (csa_tree_mul_77_11_groupi_n_299 & csa_tree_mul_77_11_groupi_n_324)));
 assign n_930 = (csa_tree_mul_77_11_groupi_n_345 ^ (csa_tree_mul_77_11_groupi_n_299 ^ csa_tree_mul_77_11_groupi_n_324));
 assign n_1352 = ((csa_tree_add_86_2_n_728 & csa_tree_add_86_2_n_721) | ((csa_tree_add_86_2_n_721 & csa_tree_add_86_2_n_637)
    | (csa_tree_add_86_2_n_637 & csa_tree_add_86_2_n_728)));
 assign n_1008 = (csa_tree_add_86_2_n_721 ^ (csa_tree_add_86_2_n_637 ^ csa_tree_add_86_2_n_728));
 assign csa_tree_mul_77_11_groupi_n_473 = ((n_348 & n_345) | ((n_345 & n_164) | (n_164 & n_348)));
 assign csa_tree_mul_77_11_groupi_n_474 = (n_345 ^ (n_164 ^ n_348));
 assign n_941 = ((csa_tree_add_106_2_groupi_n_1006 & csa_tree_add_106_2_groupi_n_957) | ((csa_tree_add_106_2_groupi_n_957
    & csa_tree_add_106_2_groupi_n_993) | (csa_tree_add_106_2_groupi_n_993 & csa_tree_add_106_2_groupi_n_1006)));
 assign n_940 = (csa_tree_add_106_2_groupi_n_957 ^ (csa_tree_add_106_2_groupi_n_993 ^ csa_tree_add_106_2_groupi_n_1006));
 assign n_998 = ((csa_tree_add_106_2_groupi_n_602 & csa_tree_add_106_2_groupi_n_762) | ((csa_tree_add_106_2_groupi_n_762
    & csa_tree_add_106_2_groupi_n_717) | (csa_tree_add_106_2_groupi_n_717 & csa_tree_add_106_2_groupi_n_602)));
 assign n_997 = (csa_tree_add_106_2_groupi_n_762 ^ (csa_tree_add_106_2_groupi_n_717 ^ csa_tree_add_106_2_groupi_n_602));
 assign n_961 = ((csa_tree_add_92_2_groupi_n_168 & csa_tree_add_92_2_groupi_n_147) | ((csa_tree_add_92_2_groupi_n_147
    & csa_tree_add_92_2_groupi_n_140) | (csa_tree_add_92_2_groupi_n_140 & csa_tree_add_92_2_groupi_n_168)));
 assign n_960 = (csa_tree_add_92_2_groupi_n_147 ^ (csa_tree_add_92_2_groupi_n_140 ^ csa_tree_add_92_2_groupi_n_168));
 assign n_1011 = ((csa_tree_add_106_2_groupi_n_683 & csa_tree_add_106_2_groupi_n_736) | ((csa_tree_add_106_2_groupi_n_736
    & csa_tree_add_106_2_groupi_n_747) | (csa_tree_add_106_2_groupi_n_747 & csa_tree_add_106_2_groupi_n_683)));
 assign n_1010 = (csa_tree_add_106_2_groupi_n_736 ^ (csa_tree_add_106_2_groupi_n_747 ^ csa_tree_add_106_2_groupi_n_683));
 assign n_962 = ((csa_tree_mul_77_11_groupi_n_395 & csa_tree_mul_77_11_groupi_n_402) | ((csa_tree_mul_77_11_groupi_n_402
    & csa_tree_mul_77_11_groupi_n_357) | (csa_tree_mul_77_11_groupi_n_357 & csa_tree_mul_77_11_groupi_n_395)));
 assign n_794 = (csa_tree_mul_77_11_groupi_n_402 ^ (csa_tree_mul_77_11_groupi_n_357 ^ csa_tree_mul_77_11_groupi_n_395));
 assign n_953 = ((csa_tree_add_92_2_groupi_n_146 & csa_tree_add_92_2_groupi_n_145) | ((csa_tree_add_92_2_groupi_n_145
    & csa_tree_add_92_2_groupi_n_120) | (csa_tree_add_92_2_groupi_n_120 & csa_tree_add_92_2_groupi_n_146)));
 assign n_952 = (csa_tree_add_92_2_groupi_n_145 ^ (csa_tree_add_92_2_groupi_n_120 ^ csa_tree_add_92_2_groupi_n_146));
 assign n_980 = ((csa_tree_add_106_2_groupi_n_630 & csa_tree_add_106_2_groupi_n_385) | ((csa_tree_add_106_2_groupi_n_385
    & csa_tree_add_106_2_groupi_n_384) | (csa_tree_add_106_2_groupi_n_384 & csa_tree_add_106_2_groupi_n_630)));
 assign n_979 = (csa_tree_add_106_2_groupi_n_385 ^ (csa_tree_add_106_2_groupi_n_384 ^ csa_tree_add_106_2_groupi_n_630));
 assign n_1000 = ((csa_tree_add_86_2_n_132 & csa_tree_add_86_2_n_156) | ((csa_tree_add_86_2_n_156 & csa_tree_add_86_2_n_874)
    | (csa_tree_add_86_2_n_874 & csa_tree_add_86_2_n_132)));
 assign n_999 = (csa_tree_add_86_2_n_156 ^ (csa_tree_add_86_2_n_874 ^ csa_tree_add_86_2_n_132));
 assign n_970 = ((csa_tree_add_92_2_groupi_n_183 & csa_tree_add_92_2_groupi_n_206) | ((csa_tree_add_92_2_groupi_n_206
    & csa_tree_add_92_2_groupi_n_186) | (csa_tree_add_92_2_groupi_n_186 & csa_tree_add_92_2_groupi_n_183)));
 assign n_969 = (csa_tree_add_92_2_groupi_n_206 ^ (csa_tree_add_92_2_groupi_n_186 ^ csa_tree_add_92_2_groupi_n_183));
 assign n_973 = ((csa_tree_add_86_2_n_643 & csa_tree_add_86_2_n_741) | ((csa_tree_add_86_2_n_741 & csa_tree_add_86_2_n_734)
    | (csa_tree_add_86_2_n_734 & csa_tree_add_86_2_n_643)));
 assign n_782 = (csa_tree_add_86_2_n_741 ^ (csa_tree_add_86_2_n_734 ^ csa_tree_add_86_2_n_643));
 assign n_990 = ((csa_tree_add_92_2_groupi_n_158 & csa_tree_add_92_2_groupi_n_169) | ((csa_tree_add_92_2_groupi_n_169
    & csa_tree_add_92_2_groupi_n_141) | (csa_tree_add_92_2_groupi_n_141 & csa_tree_add_92_2_groupi_n_158)));
 assign n_989 = (csa_tree_add_92_2_groupi_n_169 ^ (csa_tree_add_92_2_groupi_n_141 ^ csa_tree_add_92_2_groupi_n_158));
 assign n_929 = ((csa_tree_add_86_2_n_893 & csa_tree_add_86_2_n_882) | ((csa_tree_add_86_2_n_882 & csa_tree_add_86_2_n_888)
    | (csa_tree_add_86_2_n_888 & csa_tree_add_86_2_n_893)));
 assign n_928 = (csa_tree_add_86_2_n_882 ^ (csa_tree_add_86_2_n_888 ^ csa_tree_add_86_2_n_893));
 assign n_684 = ((n_1385 & final_adder_add_86_2_n_49) | ((final_adder_add_86_2_n_49 & n_1354) | (n_1354
    & n_1385)));
 assign n_717 = (final_adder_add_86_2_n_49 ^ (n_1354 ^ n_1385));
 assign n_978 = ((csa_tree_add_86_2_n_677 & csa_tree_add_86_2_n_693) | ((csa_tree_add_86_2_n_693 & csa_tree_add_86_2_n_740)
    | (csa_tree_add_86_2_n_740 & csa_tree_add_86_2_n_677)));
 assign n_977 = (csa_tree_add_86_2_n_693 ^ (csa_tree_add_86_2_n_740 ^ csa_tree_add_86_2_n_677));
 assign n_1009 = ((n_40 & n_44) | ((n_44 & n_33) | (n_33 & n_40)));
 assign n_1458 = (n_44 ^ (n_33 ^ n_40));
 assign n_939 = ((csa_tree_add_86_2_n_869 & csa_tree_add_86_2_n_895) | ((csa_tree_add_86_2_n_895 & csa_tree_add_86_2_n_884)
    | (csa_tree_add_86_2_n_884 & csa_tree_add_86_2_n_869)));
 assign n_780 = (csa_tree_add_86_2_n_895 ^ (csa_tree_add_86_2_n_884 ^ csa_tree_add_86_2_n_869));
 assign n_927 = ((csa_tree_add_86_2_n_868 & csa_tree_add_86_2_n_863) | ((csa_tree_add_86_2_n_863 & csa_tree_add_86_2_n_859)
    | (csa_tree_add_86_2_n_859 & csa_tree_add_86_2_n_868)));
 assign n_926 = (csa_tree_add_86_2_n_863 ^ (csa_tree_add_86_2_n_859 ^ csa_tree_add_86_2_n_868));
 assign n_1002 = ((csa_tree_add_86_2_n_886 & csa_tree_add_86_2_n_883) | ((csa_tree_add_86_2_n_883 & csa_tree_add_86_2_n_889)
    | (csa_tree_add_86_2_n_889 & csa_tree_add_86_2_n_886)));
 assign n_1001 = (csa_tree_add_86_2_n_883 ^ (csa_tree_add_86_2_n_889 ^ csa_tree_add_86_2_n_886));
 assign csa_tree_add_106_2_groupi_n_830 = ((csa_tree_add_106_2_groupi_n_735 & csa_tree_add_106_2_groupi_n_740)
    | ((csa_tree_add_106_2_groupi_n_740 & csa_tree_add_106_2_groupi_n_681) | (csa_tree_add_106_2_groupi_n_681
    & csa_tree_add_106_2_groupi_n_735)));
 assign n_949 = (csa_tree_add_106_2_groupi_n_740 ^ (csa_tree_add_106_2_groupi_n_681 ^ csa_tree_add_106_2_groupi_n_735));
 assign n_976 = ((csa_tree_add_86_2_n_673 & csa_tree_add_86_2_n_729) | ((csa_tree_add_86_2_n_729 & csa_tree_add_86_2_n_692)
    | (csa_tree_add_86_2_n_692 & csa_tree_add_86_2_n_673)));
 assign n_975 = (csa_tree_add_86_2_n_729 ^ (csa_tree_add_86_2_n_692 ^ csa_tree_add_86_2_n_673));
 assign n_957 = ((csa_tree_mul_77_11_groupi_n_215 & csa_tree_mul_77_11_groupi_n_205) | ((csa_tree_mul_77_11_groupi_n_205
    & csa_tree_mul_77_11_groupi_n_254) | (csa_tree_mul_77_11_groupi_n_254 & csa_tree_mul_77_11_groupi_n_215)));
 assign n_956 = (csa_tree_mul_77_11_groupi_n_205 ^ (csa_tree_mul_77_11_groupi_n_254 ^ csa_tree_mul_77_11_groupi_n_215));
 assign n_968 = ((csa_tree_add_86_2_n_830 & csa_tree_add_86_2_n_844) | ((csa_tree_add_86_2_n_844 & csa_tree_add_86_2_n_833)
    | (csa_tree_add_86_2_n_833 & csa_tree_add_86_2_n_830)));
 assign n_967 = (csa_tree_add_86_2_n_844 ^ (csa_tree_add_86_2_n_833 ^ csa_tree_add_86_2_n_830));
 assign final_adder_add_69_2_n_6 = (({in2[3]} & final_adder_add_69_2_n_4) | ((final_adder_add_69_2_n_4
    & {in1[3]}) | ({in1[3]} & {in2[3]})));
 assign n_1435 = (final_adder_add_69_2_n_4 ^ ({in1[3]} ^ {in2[3]}));
 assign n_964 = ((csa_tree_add_86_2_n_198 & csa_tree_add_86_2_n_109) | ((csa_tree_add_86_2_n_109 & csa_tree_add_86_2_n_182)
    | (csa_tree_add_86_2_n_182 & csa_tree_add_86_2_n_198)));
 assign n_963 = (csa_tree_add_86_2_n_109 ^ (csa_tree_add_86_2_n_182 ^ csa_tree_add_86_2_n_198));
 assign n_1351 = ((csa_tree_add_86_2_n_720 & csa_tree_add_86_2_n_705) | ((csa_tree_add_86_2_n_705 & csa_tree_add_86_2_n_636)
    | (csa_tree_add_86_2_n_636 & csa_tree_add_86_2_n_720)));
 assign n_1380 = (csa_tree_add_86_2_n_705 ^ (csa_tree_add_86_2_n_636 ^ csa_tree_add_86_2_n_720));
 assign n_982 = ((csa_tree_add_86_2_n_772 & csa_tree_add_86_2_n_232) | ((csa_tree_add_86_2_n_232 & csa_tree_add_86_2_n_556)
    | (csa_tree_add_86_2_n_556 & csa_tree_add_86_2_n_772)));
 assign n_981 = (csa_tree_add_86_2_n_232 ^ (csa_tree_add_86_2_n_556 ^ csa_tree_add_86_2_n_772));
 assign n_938 = ((csa_tree_add_106_2_groupi_n_687 & csa_tree_add_106_2_groupi_n_554) | ((csa_tree_add_106_2_groupi_n_554
    & csa_tree_add_106_2_groupi_n_553) | (csa_tree_add_106_2_groupi_n_553 & csa_tree_add_106_2_groupi_n_687)));
 assign n_937 = (csa_tree_add_106_2_groupi_n_554 ^ (csa_tree_add_106_2_groupi_n_553 ^ csa_tree_add_106_2_groupi_n_687));
 assign n_796 = (({in2[7]} & final_adder_add_69_2_n_12) | ((final_adder_add_69_2_n_12 & {in1[7]}) | ({in1[7]}
    & {in2[7]})));
 assign n_1431 = (final_adder_add_69_2_n_12 ^ ({in1[7]} ^ {in2[7]}));
 assign n_972 = ((csa_tree_add_106_2_groupi_n_778 & csa_tree_add_106_2_groupi_n_497) | ((csa_tree_add_106_2_groupi_n_497
    & csa_tree_add_106_2_groupi_n_771) | (csa_tree_add_106_2_groupi_n_771 & csa_tree_add_106_2_groupi_n_778)));
 assign n_971 = (csa_tree_add_106_2_groupi_n_497 ^ (csa_tree_add_106_2_groupi_n_771 ^ csa_tree_add_106_2_groupi_n_778));
 assign n_988 = ((csa_tree_add_86_2_n_862 & csa_tree_add_86_2_n_855) | ((csa_tree_add_86_2_n_855 & csa_tree_add_86_2_n_858)
    | (csa_tree_add_86_2_n_858 & csa_tree_add_86_2_n_862)));
 assign n_987 = (csa_tree_add_86_2_n_855 ^ (csa_tree_add_86_2_n_858 ^ csa_tree_add_86_2_n_862));
 assign add_100_2_n_26 = (({in4[1]} & add_100_2_n_22) | ((add_100_2_n_22 & {in3[1]}) | ({in3[1]} & {in4[1]})));
 assign n_1446 = (add_100_2_n_22 ^ ({in3[1]} ^ {in4[1]}));
 assign n_935 = ((csa_tree_mul_77_11_groupi_n_304 & csa_tree_mul_77_11_groupi_n_285) | ((csa_tree_mul_77_11_groupi_n_285
    & csa_tree_mul_77_11_groupi_n_356) | (csa_tree_mul_77_11_groupi_n_356 & csa_tree_mul_77_11_groupi_n_304)));
 assign n_934 = (csa_tree_mul_77_11_groupi_n_285 ^ (csa_tree_mul_77_11_groupi_n_356 ^ csa_tree_mul_77_11_groupi_n_304));
 assign n_966 = ((csa_tree_add_106_2_groupi_n_599 & csa_tree_add_106_2_groupi_n_437) | ((csa_tree_add_106_2_groupi_n_437
    & csa_tree_add_106_2_groupi_n_761) | (csa_tree_add_106_2_groupi_n_761 & csa_tree_add_106_2_groupi_n_599)));
 assign n_965 = (csa_tree_add_106_2_groupi_n_437 ^ (csa_tree_add_106_2_groupi_n_761 ^ csa_tree_add_106_2_groupi_n_599));
 assign n_933 = ((csa_tree_add_106_2_groupi_n_696 & csa_tree_add_106_2_groupi_n_462) | ((csa_tree_add_106_2_groupi_n_462
    & csa_tree_add_106_2_groupi_n_637) | (csa_tree_add_106_2_groupi_n_637 & csa_tree_add_106_2_groupi_n_696)));
 assign n_932 = (csa_tree_add_106_2_groupi_n_462 ^ (csa_tree_add_106_2_groupi_n_637 ^ csa_tree_add_106_2_groupi_n_696));
 assign n_1368 = ((n_121 & n_145) | ((n_145 & n_138) | (n_138 & n_121)));
 assign n_1400 = (n_145 ^ (n_138 ^ n_121));
 assign n_1005 = ((csa_tree_mul_77_11_groupi_n_212 & csa_tree_mul_77_11_groupi_n_224) | ((csa_tree_mul_77_11_groupi_n_224
    & csa_tree_mul_77_11_groupi_n_256) | (csa_tree_mul_77_11_groupi_n_256 & csa_tree_mul_77_11_groupi_n_212)));
 assign n_1004 = (csa_tree_mul_77_11_groupi_n_224 ^ (csa_tree_mul_77_11_groupi_n_256 ^ csa_tree_mul_77_11_groupi_n_212));
 assign n_1369 = ((n_436 & n_112) | ((n_112 & n_122) | (n_122 & n_436)));
 assign n_657 = (n_112 ^ (n_122 ^ n_436));
 assign final_adder_add_69_2_n_10 = (({in2[5]} & final_adder_add_69_2_n_8) | ((final_adder_add_69_2_n_8
    & {in1[5]}) | ({in1[5]} & {in2[5]})));
 assign n_1433 = (final_adder_add_69_2_n_8 ^ ({in1[5]} ^ {in2[5]}));
 assign n_1013 = ((csa_tree_add_106_2_groupi_n_967 & csa_tree_add_106_2_groupi_n_994) | ((csa_tree_add_106_2_groupi_n_994
    & csa_tree_add_106_2_groupi_n_991) | (csa_tree_add_106_2_groupi_n_991 & csa_tree_add_106_2_groupi_n_967)));
 assign n_1012 = (csa_tree_add_106_2_groupi_n_994 ^ (csa_tree_add_106_2_groupi_n_991 ^ csa_tree_add_106_2_groupi_n_967));
 assign n_944 = ((n_1377 & n_1407) | ((n_1407 & csa_tree_add_92_2_groupi_n_31) | (csa_tree_add_92_2_groupi_n_31
    & n_1377)));
 assign n_943 = (n_1407 ^ (csa_tree_add_92_2_groupi_n_31 ^ n_1377));
 assign n_992 = ((csa_tree_add_92_2_groupi_n_109 & csa_tree_add_92_2_groupi_n_144) | ((csa_tree_add_92_2_groupi_n_144
    & csa_tree_add_92_2_groupi_n_106) | (csa_tree_add_92_2_groupi_n_106 & csa_tree_add_92_2_groupi_n_109)));
 assign n_991 = (csa_tree_add_92_2_groupi_n_144 ^ (csa_tree_add_92_2_groupi_n_106 ^ csa_tree_add_92_2_groupi_n_109));
 assign n_948 = ((csa_tree_add_92_2_groupi_n_42 & csa_tree_add_92_2_groupi_n_108) | ((csa_tree_add_92_2_groupi_n_108
    & csa_tree_add_92_2_groupi_n_11) | (csa_tree_add_92_2_groupi_n_11 & csa_tree_add_92_2_groupi_n_42)));
 assign n_947 = (csa_tree_add_92_2_groupi_n_108 ^ (csa_tree_add_92_2_groupi_n_11 ^ csa_tree_add_92_2_groupi_n_42));
 assign n_996 = ((csa_tree_mul_77_11_groupi_n_192 & csa_tree_mul_77_11_groupi_n_331) | ((csa_tree_mul_77_11_groupi_n_331
    & csa_tree_mul_77_11_groupi_n_250) | (csa_tree_mul_77_11_groupi_n_250 & csa_tree_mul_77_11_groupi_n_192)));
 assign n_995 = (csa_tree_mul_77_11_groupi_n_331 ^ (csa_tree_mul_77_11_groupi_n_250 ^ csa_tree_mul_77_11_groupi_n_192));
 assign n_786 = ((n_797 & n_344) | ((n_344 & n_798) | (n_798 & n_797)));
 assign csa_tree_mul_77_11_groupi_n_457 = (n_344 ^ (n_798 ^ n_797));
 assign n_984 = ((csa_tree_add_86_2_n_819 & csa_tree_add_86_2_n_243) | ((csa_tree_add_86_2_n_243 & csa_tree_add_86_2_n_832)
    | (csa_tree_add_86_2_n_832 & csa_tree_add_86_2_n_819)));
 assign n_983 = (csa_tree_add_86_2_n_243 ^ (csa_tree_add_86_2_n_832 ^ csa_tree_add_86_2_n_819));
 assign n_955 = ((csa_tree_add_86_2_n_382 & csa_tree_add_86_2_n_174) | ((csa_tree_add_86_2_n_174 & csa_tree_add_86_2_n_250)
    | (csa_tree_add_86_2_n_250 & csa_tree_add_86_2_n_382)));
 assign n_954 = (csa_tree_add_86_2_n_174 ^ (csa_tree_add_86_2_n_250 ^ csa_tree_add_86_2_n_382));
 assign n_994 = ((csa_tree_add_86_2_n_818 & csa_tree_add_86_2_n_233) | ((csa_tree_add_86_2_n_233 & csa_tree_add_86_2_n_773)
    | (csa_tree_add_86_2_n_773 & csa_tree_add_86_2_n_818)));
 assign n_993 = (csa_tree_add_86_2_n_233 ^ (csa_tree_add_86_2_n_773 ^ csa_tree_add_86_2_n_818));
 assign mul_109_11_n_466 = ~((n_734 | n_720) & (n_732 | n_86));
 assign mul_109_11_n_477 = ~((n_728 | n_720) & (n_227 | n_86));
 assign mul_109_11_n_470 = ~((n_724 | n_720) & (n_727 | n_86));
 assign mul_109_11_n_546 = ~((n_750 | n_585) & (n_232 | n_311));
 assign n_1154 = ~(n_1156 & ~(n_1155 & csa_tree_add_92_2_groupi_n_197));
 assign mul_109_11_n_548 = ~((mul_109_11_n_383 & n_1173) | (mul_109_11_n_169 & n_370));
 assign csa_tree_add_106_2_groupi_n_374 = ~(n_803 & ~(csa_tree_add_106_2_groupi_n_69 & n_1168));
 assign csa_tree_mul_77_11_groupi_n_613 = ~(n_131 & (csa_tree_mul_77_11_groupi_n_604 | n_374));
 assign mul_109_11_n_551 = ~(n_1145 | (mul_109_11_n_41 | (mul_109_11_n_62 & n_37)));
 assign mul_109_11_n_597 = ~(n_1174 | (n_229 | (mul_109_11_n_65 & n_388)));
 assign csa_tree_add_106_2_groupi_n_372 = ~(n_1167 & ((n_233 | n_412) & (n_1118 | n_414)));
 assign mul_109_11_n_552 = ~(mul_109_11_n_43 | (n_1142 | (n_45 & mul_109_11_n_63)));
 assign csa_tree_add_106_2_groupi_n_343 = ~(csa_tree_add_106_2_groupi_n_226 & ~csa_tree_add_106_2_groupi_n_212);
 assign csa_tree_add_106_2_groupi_n_1 = ~(csa_tree_add_106_2_groupi_n_224 & ~csa_tree_add_106_2_groupi_n_220);
 assign n_1014 = ~(n_111 ^ n_1069);
 assign n_687 = ~(n_801 & ~csa_tree_add_92_2_groupi_n_81);
 assign n_1148 = ~(n_1150 & ~(n_1149 & n_118));
 assign n_1015 = ~(n_1016 ^ csa_tree_add_92_2_groupi_n_197);
 assign n_692 = ~(csa_tree_add_92_2_groupi_n_82 ^ n_802);
 assign n_1147 = ~(n_1150 & ~(n_111 & n_1149));
 assign n_1427 = ~(n_1069 ^ n_118);
 assign n_716 = ~(n_852 ^ n_68);
 assign mul_109_11_n_476 = ~((n_585 | n_767) & (n_763 | n_311));
 assign mul_109_11_n_463 = ~((n_720 | n_721) & (n_722 | n_86));
 assign mul_109_11_n_462 = ~((n_720 | n_722) & (n_729 | n_86));
 assign mul_109_11_n_461 = ~((n_720 | n_738) & (n_735 | n_86));
 assign mul_109_11_n_460 = ~((n_730 | n_720) & (n_725 | n_86));
 assign mul_109_11_n_459 = ~((n_726 | n_720) & (n_723 | n_86));
 assign mul_109_11_n_458 = ~((n_723 | n_720) & (n_724 | n_86));
 assign mul_109_11_n_457 = ~((n_725 | n_720) & (n_726 | n_86));
 assign mul_109_11_n_456 = ~((n_742 | n_720) & (n_737 | n_86));
 assign mul_109_11_n_454 = ~((n_235 | n_720) & (n_733 | n_86));
 assign mul_109_11_n_453 = ~((n_727 | n_720) & (n_728 | n_86));
 assign mul_109_11_n_452 = ~((n_720 | n_731) & (n_741 | n_86));
 assign mul_109_11_n_451 = ~((n_720 | n_729) & (n_730 | n_86));
 assign mul_109_11_n_450 = ~((n_720 | n_740) & (n_731 | n_86));
 assign mul_109_11_n_445 = ~((n_732 | n_720) & (n_739 | n_86));
 assign mul_109_11_n_443 = ~((n_733 | n_720) & (n_734 | n_86));
 assign mul_109_11_n_440 = ~((n_720 | n_737) & (n_738 | n_86));
 assign mul_109_11_n_442 = ~((n_720 | n_735) & (n_736 | n_86));
 assign mul_109_11_n_439 = ~((n_720 | n_739) & (n_740 | n_86));
 assign mul_109_11_n_434 = ~((n_720 | n_741) & (n_742 | n_86));
 assign mul_109_11_n_519 = ~((n_759 | n_585) & (n_719 | n_311));
 assign mul_109_11_n_480 = ~((n_752 | n_585) & (n_773 | n_311));
 assign mul_109_11_n_478 = ~((n_228 | n_585) & (n_752 | n_311));
 assign mul_109_11_n_464 = ~((n_720 | n_736) & (n_721 | n_86));
 assign mul_109_11_n_474 = ~((n_764 | n_585) & (n_753 | n_311));
 assign mul_109_11_n_473 = ~((n_585 | n_753) & (n_760 | n_311));
 assign mul_109_11_n_472 = ~((n_585 | n_756) & (n_771 | n_311));
 assign mul_109_11_n_471 = ~((n_585 | n_754) & (n_755 | n_311));
 assign mul_109_11_n_467 = ~((n_585 | n_768) & (n_766 | n_311));
 assign mul_109_11_n_455 = ~((n_585 | n_758) & (n_754 | n_311));
 assign mul_109_11_n_438 = ~((n_585 | n_755) & (n_775 | n_311));
 assign mul_109_11_n_435 = ~((n_757 | n_585) & (n_769 | n_311));
 assign mul_109_11_n_433 = ~((n_762 | n_585) & (n_756 | n_311));
 assign mul_109_11_n_432 = ~((n_772 | n_585) & (n_757 | n_311));
 assign mul_109_11_n_430 = ~((n_585 | n_761) & (n_758 | n_311));
 assign mul_109_11_n_429 = ~((n_765 | n_585) & (n_759 | n_311));
 assign mul_109_11_n_428 = ~((n_585 | n_760) & (n_761 | n_311));
 assign mul_109_11_n_427 = ~((n_585 | n_776) & (n_762 | n_311));
 assign mul_109_11_n_424 = ~((n_585 | n_763) & (n_764 | n_311));
 assign mul_109_11_n_422 = ~((n_770 | n_585) & (n_765 | n_311));
 assign mul_109_11_n_421 = ~((n_585 | n_766) & (n_767 | n_311));
 assign mul_109_11_n_419 = ~((n_774 | n_585) & (n_768 | n_311));
 assign mul_109_11_n_418 = ~((n_769 | n_585) & (n_770 | n_311));
 assign mul_109_11_n_417 = ~((n_585 | n_771) & (n_772 | n_311));
 assign mul_109_11_n_415 = ~((n_773 | n_585) & (n_774 | n_311));
 assign mul_109_11_n_414 = ~((n_585 | n_775) & (n_776 | n_311));
 assign mul_109_11_n_550 = ~(n_1185 | ((n_362 & n_201) | (mul_109_11_n_61 & n_84)));
 assign csa_tree_add_106_2_groupi_n_516 = ~((n_877 | n_371) & (n_874 | n_435));
 assign csa_tree_add_106_2_groupi_n_551 = ~((n_893 | n_399) & (n_898 | n_397));
 assign csa_tree_add_106_2_groupi_n_550 = ~((n_1102 | n_399) & (n_1105 | n_397));
 assign csa_tree_add_106_2_groupi_n_549 = ~((n_1101 | n_399) & (n_1102 | n_397));
 assign csa_tree_add_106_2_groupi_n_546 = ~((n_1104 | n_399) & (n_1100 | n_397));
 assign csa_tree_add_106_2_groupi_n_543 = ~((n_1103 | n_397) & (n_1100 | n_399));
 assign csa_tree_add_106_2_groupi_n_527 = ~((n_1098 | n_391) & (n_1099 | n_389));
 assign csa_tree_add_106_2_groupi_n_517 = ~((n_1095 | n_391) & (n_1096 | n_389));
 assign csa_tree_add_106_2_groupi_n_512 = ~((n_891 | n_389) & (n_892 | n_391));
 assign csa_tree_add_106_2_groupi_n_507 = ~((n_1095 | n_389) & (n_1094 | n_391));
 assign csa_tree_add_106_2_groupi_n_506 = ~((n_890 | n_391) & (n_892 | n_389));
 assign csa_tree_add_106_2_groupi_n_502 = ~((n_1093 | n_389) & (n_1099 | n_391));
 assign csa_tree_add_106_2_groupi_n_492 = ~((n_1091 | n_389) & (n_1090 | n_391));
 assign csa_tree_add_106_2_groupi_n_490 = ~((n_1092 | n_391) & (n_1094 | n_389));
 assign csa_tree_add_106_2_groupi_n_489 = ~((n_888 | n_391) & (n_889 | n_389));
 assign csa_tree_add_106_2_groupi_n_488 = ~((n_1091 | n_391) & (n_1092 | n_389));
 assign csa_tree_add_106_2_groupi_n_484 = ~((n_1093 | n_391) & (n_1090 | n_389));
 assign csa_tree_add_106_2_groupi_n_458 = ~((n_1088 | n_380) & (n_1089 | n_378));
 assign csa_tree_mul_77_11_groupi_n_601 = (n_248 | (csa_tree_mul_77_11_groupi_n_590 & csa_tree_mul_77_11_groupi_n_522));
 assign mul_109_11_n_666 = ~(n_1162 | n_1175);
 assign mul_109_11_n_672 = ~(n_1017 | n_1176);
 assign mul_109_11_n_664 = (n_82 & (n_1169 | n_1034));
 assign mul_109_11_n_395 = ~(n_1160 | mul_109_11_n_39);
 assign mul_109_11_n_665 = ~(n_1152 | n_1183);
 assign mul_109_11_n_671 = ~(n_1161 | mul_109_11_n_25);
 assign n_801 = ~(n_802 & (n_51 | n_10));
 assign csa_tree_add_106_2_groupi_n_457 = ~((n_1086 | n_380) & (n_1087 | n_378));
 assign csa_tree_add_106_2_groupi_n_5 = ((n_1124 | n_427) & (n_259 | n_441));
 assign csa_tree_add_106_2_groupi_n_454 = ~((n_1088 | n_378) & (n_1085 | n_380));
 assign csa_tree_add_106_2_groupi_n_500 = ~((n_889 | n_391) & (n_890 | n_389));
 assign csa_tree_add_106_2_groupi_n_453 = ~((n_1040 | n_378) & (n_1121 | n_380));
 assign csa_tree_add_106_2_groupi_n_452 = ~((n_886 | n_378) & (n_887 | n_380));
 assign n_803 = ~((n_1412 & (n_1470 & n_418)) | (n_1323 & n_1478));
 assign csa_tree_add_106_2_groupi_n_450 = ~((n_884 | n_380) & (n_885 | n_378));
 assign csa_tree_add_106_2_groupi_n_449 = ~((n_1083 | n_380) & (n_1084 | n_378));
 assign csa_tree_add_106_2_groupi_n_448 = ~((n_1120 | n_380) & (n_1121 | n_378));
 assign csa_tree_add_106_2_groupi_n_447 = ~((n_1087 | n_380) & (n_1082 | n_378));
 assign csa_tree_add_106_2_groupi_n_443 = ~((n_1061 | n_380) & (n_1120 | n_378));
 assign csa_tree_add_106_2_groupi_n_442 = ~((n_885 | n_380) & (n_887 | n_378));
 assign csa_tree_add_106_2_groupi_n_441 = ~((n_1061 | n_378) & (n_1082 | n_380));
 assign csa_tree_add_106_2_groupi_n_569 = ~((n_1106 | n_399) & (n_1107 | n_397));
 assign csa_tree_add_106_2_groupi_n_440 = ~((n_1086 | n_378) & (n_1089 | n_380));
 assign csa_tree_add_106_2_groupi_n_435 = ~((n_1084 | n_380) & (n_1085 | n_378));
 assign csa_tree_add_106_2_groupi_n_524 = ~((n_1097 | n_391) & (n_1098 | n_389));
 assign csa_tree_add_106_2_groupi_n_609 = ~((n_1079 | n_371) & (n_1080 | n_435));
 assign csa_tree_add_106_2_groupi_n_626 = ~((n_1079 | n_435) & (n_234 | n_371));
 assign csa_tree_add_106_2_groupi_n_535 = ~((n_882 | n_371) & (n_883 | n_435));
 assign csa_tree_add_106_2_groupi_n_533 = ~((n_1077 | n_435) & (n_1078 | n_371));
 assign csa_tree_add_106_2_groupi_n_532 = ~((n_880 | n_435) & (n_883 | n_371));
 assign csa_tree_add_106_2_groupi_n_486 = ~((n_872 | n_435) & (n_873 | n_371));
 assign csa_tree_add_106_2_groupi_n_494 = ~((n_873 | n_435) & (n_874 | n_371));
 assign csa_tree_add_106_2_groupi_n_495 = ~((n_1072 | n_435) & (n_1075 | n_371));
 assign csa_tree_add_106_2_groupi_n_501 = ~((n_1070 | n_435) & (n_1071 | n_371));
 assign csa_tree_add_106_2_groupi_n_508 = ~((n_1071 | n_435) & (n_1072 | n_371));
 assign csa_tree_add_106_2_groupi_n_510 = ~((n_875 | n_371) & (n_876 | n_435));
 assign csa_tree_add_106_2_groupi_n_511 = ~((n_879 | n_371) & (n_877 | n_435));
 assign csa_tree_add_106_2_groupi_n_513 = ~((n_1076 | n_435) & (n_1080 | n_371));
 assign csa_tree_add_106_2_groupi_n_514 = ~((n_881 | n_371) & (n_878 | n_435));
 assign csa_tree_add_106_2_groupi_n_531 = ~((n_1078 | n_435) & (n_1076 | n_371));
 assign csa_tree_add_106_2_groupi_n_520 = ~((n_879 | n_435) & (n_1074 | n_371));
 assign csa_tree_add_106_2_groupi_n_523 = ~((n_880 | n_371) & (n_881 | n_435));
 assign csa_tree_add_106_2_groupi_n_526 = ~((n_1073 | n_371) & (n_1074 | n_435));
 assign csa_tree_add_106_2_groupi_n_528 = ~((n_1077 | n_371) & (n_1075 | n_435));
 assign csa_tree_add_106_2_groupi_n_529 = ~((n_882 | n_435) & (n_872 | n_371));
 assign csa_tree_add_106_2_groupi_n_530 = ~((n_1070 | n_371) & (n_1073 | n_435));
 assign csa_tree_add_106_2_groupi_n_119 = ~((n_1347 | n_1440) & (csa_tree_add_106_2_groupi_n_48 | csa_tree_add_106_2_groupi_n_43));
 assign csa_tree_add_106_2_groupi_n_228 = ~(csa_tree_add_106_2_groupi_n_338 & (n_1440 | n_1439));
 assign csa_tree_add_106_2_groupi_n_94 = ~((n_1347 | n_1444) & (csa_tree_add_106_2_groupi_n_48 | csa_tree_add_106_2_groupi_n_41));
 assign csa_tree_add_106_2_groupi_n_170 = ~((n_1347 | n_1442) & (csa_tree_add_106_2_groupi_n_48 | csa_tree_add_106_2_groupi_n_42));
 assign n_715 = ~(n_851 ^ n_421);
 assign n_1018 = ~((n_1033 | n_380) & (n_1059 | n_378));
 assign n_1019 = ~((n_1096 | n_391) & (n_1044 | n_389));
 assign n_805 = ~((n_888 | n_389) & (n_391 | n_320));
 assign n_1020 = ~((n_1047 | n_399) & (n_1024 | n_397));
 assign n_806 = ~((n_841 | n_379) & (n_381 | n_65));
 assign n_1022 = ~((n_1046 | n_397) & (n_1029 | n_399));
 assign n_807 = ~((n_843 | n_423) & (n_400 | n_424));
 assign n_1023 = ~((n_1024 | n_399) & (n_1025 | n_397));
 assign n_808 = ~((n_811 | n_414) & (n_809 | n_412));
 assign n_1026 = ~((n_1031 | n_399) & (n_1028 | n_397));
 assign n_1027 = ~((n_1028 | n_399) & (n_1029 | n_397));
 assign n_810 = ~((n_811 | n_412) & (n_372 | n_414));
 assign n_1030 = ~((n_1031 | n_397) & (n_1107 | n_399));
 assign n_812 = ~((n_845 | n_378) & (n_380 | n_319));
 assign n_1032 = ~((n_1040 | n_380) & (n_1033 | n_378));
 assign n_813 = ~((n_838 | n_390) & (n_392 | n_66));
 assign n_814 = ~((n_906 | n_423) & (n_850 | n_424));
 assign n_816 = ~((n_834 | n_78) & (n_429 | n_360));
 assign csa_tree_add_106_2_groupi_n_226 = ~(n_1441 ^ n_1442);
 assign n_1041 = ~((n_247 | n_414) & (n_1042 | n_412));
 assign n_831 = ~((n_832 | n_78) & (n_835 | n_429));
 assign n_799 = ~((n_809 | n_414) & (n_901 | n_412));
 assign n_1043 = ~((n_1063 | n_389) & (n_1044 | n_391));
 assign n_1045 = ~((n_1046 | n_399) & (n_1047 | n_397));
 assign n_833 = ~((n_834 | n_429) & (n_835 | n_78));
 assign n_836 = ~((n_837 | n_390) & (n_838 | n_392));
 assign n_839 = ~((n_840 | n_379) & (n_841 | n_381));
 assign n_842 = ~((n_849 | n_423) & (n_843 | n_424));
 assign n_844 = ~((n_845 | n_380) & (n_884 | n_378));
 assign csa_tree_add_106_2_groupi_n_555 = ~((n_893 | n_397) & (n_1066 | n_399));
 assign csa_tree_add_106_2_groupi_n_587 = ~((n_1067 | n_429) & (n_821 | n_78));
 assign mul_109_11_n_612 = ~((n_870 | n_800) & (mul_109_11_n_404 | n_871));
 assign csa_tree_add_106_2_groupi_n_559 = ~((n_1103 | n_399) & (n_1106 | n_397));
 assign csa_tree_add_106_2_groupi_n_562 = ~((n_1104 | n_397) & (n_1105 | n_399));
 assign csa_tree_add_106_2_groupi_n_565 = ~((n_898 | n_399) & (n_899 | n_397));
 assign csa_tree_add_106_2_groupi_n_376 = ~((n_1109 | n_414) & (n_1110 | n_412));
 assign csa_tree_add_106_2_groupi_n_566 = ~((n_899 | n_399) & (n_897 | n_397));
 assign csa_tree_add_106_2_groupi_n_567 = ~((n_896 | n_397) & (n_897 | n_399));
 assign n_1050 = ~((n_1064 | n_391) & (n_1052 | n_389));
 assign n_1051 = ~((n_1052 | n_391) & (n_1053 | n_389));
 assign mul_109_11_n_613 = ~((mul_109_11_n_404 | n_868) & (n_869 | n_800));
 assign csa_tree_add_106_2_groupi_n_382 = ~((n_1112 | n_412) & (n_1110 | n_414));
 assign csa_tree_add_106_2_groupi_n_381 = ~((n_900 | n_412) & (n_902 | n_414));
 assign csa_tree_add_106_2_groupi_n_383 = ~((n_1113 | n_414) & (n_1119 | n_412));
 assign csa_tree_add_106_2_groupi_n_380 = ~((n_901 | n_414) & (n_902 | n_412));
 assign csa_tree_add_106_2_groupi_n_378 = ~((n_1108 | n_414) & (n_1109 | n_412));
 assign csa_tree_add_106_2_groupi_n_377 = ~((n_1108 | n_412) & (n_1111 | n_414));
 assign csa_tree_add_106_2_groupi_n_375 = ~((n_1116 | n_414) & (n_1111 | n_412));
 assign csa_tree_add_106_2_groupi_n_373 = ~((n_1112 | n_414) & (n_1113 | n_412));
 assign csa_tree_add_106_2_groupi_n_371 = ~((n_1115 | n_414) & (n_1117 | n_412));
 assign csa_tree_add_106_2_groupi_n_368 = ~((n_1114 | n_414) & (n_1115 | n_412));
 assign csa_tree_add_106_2_groupi_n_366 = ~((n_1116 | n_412) & (n_1117 | n_414));
 assign csa_tree_add_106_2_groupi_n_365 = ~((n_1118 | n_412) & (n_1119 | n_414));
 assign csa_tree_add_106_2_groupi_n_608 = ~((n_1067 | n_78) & (n_1068 | n_429));
 assign csa_tree_add_106_2_groupi_n_460 = ~((n_1129 | n_424) & (n_1130 | n_423));
 assign csa_tree_add_106_2_groupi_n_461 = ~((n_911 | n_424) & (n_905 | n_423));
 assign csa_tree_add_106_2_groupi_n_464 = ~((n_903 | n_423) & (n_904 | n_424));
 assign csa_tree_add_106_2_groupi_n_467 = ~((n_1125 | n_424) & (n_1122 | n_423));
 assign csa_tree_add_106_2_groupi_n_468 = ~((n_903 | n_424) & (n_1127 | n_423));
 assign csa_tree_add_106_2_groupi_n_470 = ~((n_1123 | n_424) & (n_1133 | n_423));
 assign csa_tree_add_106_2_groupi_n_612 = ~((n_1056 | n_78) & (n_1057 | n_429));
 assign csa_tree_add_106_2_groupi_n_471 = ~((n_1125 | n_423) & (n_1131 | n_424));
 assign csa_tree_add_106_2_groupi_n_472 = ~((n_1126 | n_423) & (n_1127 | n_424));
 assign csa_tree_add_106_2_groupi_n_475 = ~((n_904 | n_423) & (n_905 | n_424));
 assign csa_tree_add_106_2_groupi_n_476 = ~((n_907 | n_423) & (n_906 | n_424));
 assign csa_tree_add_106_2_groupi_n_477 = ~((n_907 | n_424) & (n_908 | n_423));
 assign csa_tree_add_106_2_groupi_n_478 = ~((n_909 | n_423) & (n_908 | n_424));
 assign csa_tree_add_106_2_groupi_n_479 = ~((n_1128 | n_423) & (n_1126 | n_424));
 assign csa_tree_add_106_2_groupi_n_480 = ~((n_1128 | n_424) & (n_1129 | n_423));
 assign csa_tree_add_106_2_groupi_n_481 = ~((n_909 | n_424) & (n_910 | n_423));
 assign mul_109_11_n_611 = ~((n_866 | n_800) & (mul_109_11_n_404 | n_867));
 assign csa_tree_add_106_2_groupi_n_482 = ~((n_910 | n_424) & (n_911 | n_423));
 assign csa_tree_add_106_2_groupi_n_483 = ~((n_1122 | n_424) & (n_1123 | n_423));
 assign csa_tree_add_106_2_groupi_n_485 = ~((n_1130 | n_424) & (n_1131 | n_423));
 assign csa_tree_add_106_2_groupi_n_601 = ~((n_825 | n_429) & (n_1057 | n_78));
 assign csa_tree_add_106_2_groupi_n_600 = ~((n_1038 | n_429) & (n_1039 | n_78));
 assign csa_tree_add_106_2_groupi_n_610 = ~((n_1132 | n_423) & (n_1133 | n_424));
 assign csa_tree_add_106_2_groupi_n_624 = ~((n_1138 | n_440) & (n_1134 | n_427));
 assign csa_tree_add_106_2_groupi_n_625 = ~((n_1135 | n_427) & (n_1140 | n_440));
 assign csa_tree_add_106_2_groupi_n_623 = ~((n_1136 | n_427) & (n_1135 | n_440));
 assign csa_tree_add_106_2_groupi_n_596 = ~((n_1036 | n_429) & (n_1037 | n_78));
 assign csa_tree_add_106_2_groupi_n_622 = ~((n_918 | n_427) & (n_913 | n_440));
 assign csa_tree_add_106_2_groupi_n_621 = ~((n_1137 | n_427) & (n_1136 | n_440));
 assign csa_tree_add_106_2_groupi_n_620 = ~((n_913 | n_427) & (n_914 | n_440));
 assign csa_tree_add_106_2_groupi_n_619 = ~((n_914 | n_427) & (n_915 | n_440));
 assign csa_tree_add_106_2_groupi_n_618 = ~((n_1139 | n_427) & (n_1081 | n_440));
 assign csa_tree_add_106_2_groupi_n_616 = ~((n_916 | n_440) & (n_915 | n_427));
 assign csa_tree_add_106_2_groupi_n_615 = ~((n_917 | n_440) & (n_920 | n_427));
 assign csa_tree_add_106_2_groupi_n_590 = ~((n_824 | n_78) & (n_832 | n_429));
 assign csa_tree_add_106_2_groupi_n_614 = ~((n_921 | n_440) & (n_916 | n_427));
 assign csa_tree_add_106_2_groupi_n_613 = ~((n_917 | n_427) & (n_919 | n_440));
 assign csa_tree_add_106_2_groupi_n_589 = ~((n_1048 | n_429) & (n_1049 | n_78));
 assign csa_tree_add_106_2_groupi_n_607 = ~((n_1137 | n_440) & (n_1138 | n_427));
 assign csa_tree_add_106_2_groupi_n_604 = ~((n_918 | n_440) & (n_919 | n_427));
 assign csa_tree_add_106_2_groupi_n_581 = ~((n_920 | n_440) & (n_922 | n_427));
 assign mul_109_11_n_610 = ~((n_864 | n_800) & (mul_109_11_n_404 | n_865));
 assign csa_tree_add_106_2_groupi_n_579 = ~((n_921 | n_427) & (n_1134 | n_440));
 assign csa_tree_add_106_2_groupi_n_577 = ~((n_923 | n_427) & (n_922 | n_440));
 assign csa_tree_add_106_2_groupi_n_575 = ~((n_1081 | n_427) & (n_1124 | n_440));
 assign csa_tree_add_106_2_groupi_n_572 = ~((n_1139 | n_440) & (n_1140 | n_427));
 assign mul_109_11_n_609 = ~((n_871 | n_800) & (mul_109_11_n_404 | n_863));
 assign csa_tree_add_106_2_groupi_n_570 = ~((n_923 | n_440) & (n_924 | n_427));
 assign csa_tree_add_106_2_groupi_n_588 = ~((n_822 | n_429) & (n_823 | n_78));
 assign csa_tree_add_106_2_groupi_n_585 = ~((n_1037 | n_429) & (n_1035 | n_78));
 assign csa_tree_add_106_2_groupi_n_582 = ~((n_1035 | n_429) & (n_1068 | n_78));
 assign csa_tree_add_106_2_groupi_n_574 = ~((n_822 | n_78) & (n_820 | n_429));
 assign csa_tree_add_106_2_groupi_n_571 = ~((n_1049 | n_429) & (n_1038 | n_78));
 assign csa_tree_add_106_2_groupi_n_568 = ~((n_823 | n_429) & (n_819 | n_78));
 assign csa_tree_add_106_2_groupi_n_564 = ~((n_1048 | n_78) & (n_1056 | n_429));
 assign csa_tree_add_106_2_groupi_n_556 = ~((n_824 | n_429) & (n_820 | n_78));
 assign mul_109_11_n_608 = ~((n_863 | n_800) & (mul_109_11_n_404 | n_862));
 assign csa_tree_add_106_2_groupi_n_547 = ~((n_1036 | n_78) & (n_1039 | n_429));
 assign csa_tree_add_106_2_groupi_n_544 = ~((n_817 | n_78) & (n_818 | n_429));
 assign mul_109_11_n_607 = ~((n_860 | n_800) & (mul_109_11_n_404 | n_861));
 assign csa_tree_add_106_2_groupi_n_542 = ~((n_825 | n_78) & (n_817 | n_429));
 assign csa_tree_add_106_2_groupi_n_540 = ~((n_819 | n_429) & (n_818 | n_78));
 assign mul_109_11_n_605 = ~((n_858 | n_800) & (mul_109_11_n_404 | n_859));
 assign n_1054 = ~((n_253 & n_465) | (n_265 & stall));
 assign n_1055 = ~((n_257 & n_465) | (n_1473 & stall));
 assign mul_109_11_n_595 = ~((mul_109_11_n_404 | n_857) & (n_865 | n_800));
 assign csa_tree_add_106_2_groupi_n_606 = ~((n_1132 | n_424) & (n_1494 | n_423));
 assign mul_109_11_n_593 = ~((mul_109_11_n_404 | n_860) & (n_857 | n_800));
 assign mul_109_11_n_589 = ~((n_855 | n_800) & (mul_109_11_n_404 | n_895));
 assign mul_109_11_n_554 = ~((mul_109_11_n_364 | n_800) & (mul_109_11_n_404 | n_815));
 assign mul_109_11_n_557 = ~((n_859 | n_800) & (mul_109_11_n_404 | n_870));
 assign mul_109_11_n_562 = ~((n_868 | n_800) & (mul_109_11_n_404 | n_858));
 assign mul_109_11_n_568 = ~((n_856 | n_800) & (mul_109_11_n_404 | n_864));
 assign mul_109_11_n_581 = ~((mul_109_11_n_404 | n_869) & (n_861 | n_800));
 assign mul_109_11_n_583 = ~((n_815 | n_800) & (mul_109_11_n_404 | n_854));
 assign mul_109_11_n_584 = ~((mul_109_11_n_404 | n_804) & (n_853 | n_800));
 assign mul_109_11_n_585 = ~((n_804 | n_800) & (mul_109_11_n_404 | n_230));
 assign mul_109_11_n_586 = ~((mul_109_11_n_404 | n_894) & (n_895 | n_800));
 assign mul_109_11_n_587 = ~((n_894 | n_800) & (mul_109_11_n_404 | n_853));
 assign mul_109_11_n_588 = ~((n_854 | n_800) & (mul_109_11_n_404 | n_866));
 assign mul_109_11_n_590 = ~((n_862 | n_800) & (mul_109_11_n_404 | n_855));
 assign mul_109_11_n_591 = ~((n_867 | n_800) & (mul_109_11_n_404 | n_856));
 assign n_712 = ~((n_851 | n_104) & (n_1153 | n_439));
 assign csa_tree_add_106_2_groupi_n_224 = ~(csa_tree_add_106_2_groupi_n_35 ^ csa_tree_add_106_2_groupi_n_41);
 assign n_848 = ~((n_849 | n_424) & (n_850 | n_423));
 assign n_847 = ~((n_876 | n_371) & (n_435 | n_366));
 assign n_1058 = ~((n_1059 | n_380) & (n_1060 | n_378));
 assign n_846 = ~((n_924 | n_440) & (n_427 | n_326));
 assign n_829 = ~((n_830 | n_413) & (n_415 | n_72));
 assign n_827 = ~((n_828 | n_413) & (n_830 | n_415));
 assign n_826 = ~((n_875 | n_435) & (n_878 | n_371));
 assign n_1062 = ~((n_1063 | n_391) & (n_1064 | n_389));
 assign n_1065 = ~((n_1066 | n_397) & (n_399 | n_312));
 assign mul_109_11_n_77 = ~n_1144;
 assign n_1438 = ~csa_tree_add_106_2_groupi_n_45;
 assign mul_109_11_n_79 = ~n_1141;
 assign csa_tree_add_92_2_groupi_n_81 = (n_51 & n_10);
 assign csa_tree_add_92_2_groupi_n_82 = (n_51 ^ n_10);
 assign csa_tree_add_92_2_groupi_n_91 = (n_70 & n_52);
 assign n_852 = (n_70 ^ n_52);
 assign n_1145 = (n_362 & n_1146);
 assign n_1144 = (n_362 ^ n_1146);
 assign n_1174 = (n_310 & n_362);
 assign n_1173 = (n_310 ^ n_362);
 assign n_1172 = (csa_tree_add_106_2_groupi_n_76 & csa_tree_add_106_2_groupi_n_77);
 assign n_1171 = (csa_tree_add_106_2_groupi_n_76 ^ csa_tree_add_106_2_groupi_n_77);
 assign csa_tree_add_92_2_groupi_n_89 = (n_9 & n_5);
 assign csa_tree_add_92_2_groupi_n_90 = (n_9 ^ n_5);
 assign n_1142 = (n_362 & n_1143);
 assign n_1141 = (n_362 ^ n_1143);
 assign n_1021 = ~n_1164;
 assign n_248 = ~(n_444 & (csa_tree_mul_77_11_groupi_n_537 & (n_341 | n_340)));
 assign csa_tree_mul_77_11_groupi_n_575 = ~(n_151 & (csa_tree_mul_77_11_groupi_n_572 & (n_264 | n_131)));
 assign n_226 = ~(n_1467 & (csa_tree_mul_77_11_groupi_n_368 | (csa_tree_mul_77_11_groupi_n_329 | stall)));
 assign n_216 = ~((csa_tree_mul_77_11_groupi_n_368 & (csa_tree_mul_77_11_groupi_n_329 & n_465)) | (n_252
    & stall));
 assign n_1164 = ~((n_465 & ({in8[7]} & {in7[7]})) | (n_408 & stall));
 assign n_221 = ~(n_1461 & (csa_tree_mul_77_11_groupi_n_453 | (csa_tree_mul_77_11_groupi_n_475 | stall)));
 assign n_1159 = ~(n_255 & ~(n_339 & stall));
 assign csa_tree_add_86_2_n_302 = ~(n_1153 | ~n_2);
 assign n_1165 = ~(n_1166 & n_310);
 assign n_1151 = (n_1166 | n_310);
 assign n_1160 = ~((mul_109_11_n_38 & n_1460) | (n_225 & n_1195));
 assign csa_tree_add_86_2_n_295 = ~(n_1153 | ~n_406);
 assign csa_tree_add_86_2_n_339 = ~(n_1153 | ~n_425);
 assign n_1161 = ~(n_1203 | (n_1204 & n_1199));
 assign csa_tree_add_86_2_n_289 = ~(n_1153 | ~n_430);
 assign csa_tree_mul_77_11_groupi_n_600 = ~(csa_tree_mul_77_11_groupi_n_521 & n_925);
 assign n_1152 = ~(n_1208 | (n_1209 & n_1177));
 assign mul_109_11_n_662 = ~(mul_109_11_n_56 | ((n_1451 & n_1452) | (mul_109_11_n_3 & n_362)));
 assign mul_109_11_n_661 = ~(mul_109_11_n_52 | ((mul_109_11_n_1 & n_362) | (n_1453 & n_1454)));
 assign n_1162 = ~(n_1205 | (mul_109_11_n_38 & n_1206));
 assign n_1017 = ~(n_219 | (mul_109_11_n_38 & n_1163));
 assign csa_tree_mul_77_11_groupi_n_604 = ~(csa_tree_mul_77_11_groupi_n_560 | n_925);
 assign csa_tree_add_106_2_groupi_n_338 = ~(n_1440 & n_1439);
 assign n_802 = ~(n_254 & ~(n_68 & n_52));
 assign n_720 = (n_224 | n_1474);
 assign n_585 = (n_231 | n_1472);
 assign csa_tree_add_86_2_n_7 = ~n_1341;
 assign csa_tree_add_106_2_groupi_n_41 = ~n_1444;
 assign csa_tree_add_106_2_groupi_n_43 = ~n_1440;
 assign csa_tree_add_106_2_groupi_n_42 = ~n_1442;
 assign n_851 = ~n_1153;
 assign mul_109_11_n_294 = ~((n_31 | n_310) & (n_1196 | mul_109_11_n_19));
 assign mul_109_11_n_257 = ~(n_1206 & ~n_1205);
 assign mul_109_11_n_252 = ~(n_1163 & n_220);
 assign csa_tree_mul_77_11_groupi_n_603 = ~(n_1170 & n_137);
 assign n_1167 = ~(csa_tree_add_106_2_groupi_n_68 & n_1168);
 assign mul_109_11_n_76 = ~(n_1204 & ~n_1203);
 assign mul_109_11_n_72 = ~(n_1209 & ~n_1208);
 assign mul_109_11_n_69 = ~(n_217 & ~n_1034);
 assign n_253 = ~(csa_tree_mul_77_11_groupi_n_591 & (csa_tree_mul_77_11_groupi_n_564 | csa_tree_mul_77_11_groupi_n_573));
 assign n_254 = ~(n_70 & (n_68 | n_52));
 assign n_255 = ~(n_465 & (csa_tree_mul_77_11_groupi_n_407 | csa_tree_mul_77_11_groupi_n_369));
 assign mul_109_11_n_227 = ~(n_1381 & (mul_109_11_n_56 | mul_109_11_n_38));
 assign n_1323 = ~(n_233 & ~(csa_tree_add_106_2_groupi_n_68 & n_416));
 assign csa_tree_add_106_2_groupi_n_632 = ~(n_437 & (n_429 | n_243));
 assign n_256 = ~(csa_tree_mul_77_11_groupi_n_547 ^ csa_tree_mul_77_11_groupi_n_593);
 assign n_249 = ~(csa_tree_mul_77_11_groupi_n_587 ^ csa_tree_mul_77_11_groupi_n_555);
 assign n_257 = ~(csa_tree_mul_77_11_groupi_n_328 ^ csa_tree_mul_77_11_groupi_n_174);
 assign n_258 = ~(csa_tree_add_92_2_groupi_n_32 ^ csa_tree_add_92_2_groupi_n_66);
 assign n_247 = ~((csa_tree_add_106_2_groupi_n_69 & n_416) | (n_1412 & n_418));
 assign n_246 = ~(n_387 ^ n_171);
 assign csa_tree_add_106_2_groupi_n_926 = (csa_tree_add_106_2_groupi_n_854 ^ n_62);
 assign n_245 = ~(csa_tree_add_106_2_groupi_n_767 ^ csa_tree_add_106_2_groupi_n_716);
 assign n_1169 = ~(n_218 | n_87);
 assign csa_tree_add_106_2_groupi_n_422 = ~((n_1178 | n_318) & (n_1179 | n_1182));
 assign mul_109_11_n_232 = ~((n_106 & ~n_1448) | (n_749 & n_1448));
 assign mul_109_11_n_260 = ~(n_45 ^ n_1143);
 assign csa_tree_add_106_2_groupi_n_387 = ~((csa_tree_add_106_2_groupi_n_53 | n_1179) & (n_215 | n_1178));
 assign csa_tree_add_106_2_groupi_n_408 = ~((n_202 | n_209) & (n_203 | n_210));
 assign mul_109_11_n_240 = ~((n_1146 | n_34) & (mul_109_11_n_25 | n_1199));
 assign mul_109_11_n_259 = ((mul_109_11_n_25 & ~n_37) | (n_1146 & n_37));
 assign mul_109_11_n_241 = ~((n_60 & ~n_61) | (n_1175 & n_61));
 assign mul_109_11_n_258 = ~((n_34 | n_60) & (n_1199 | n_1175));
 assign mul_109_11_n_0 = ~((n_362 & ~n_1448) | (mul_109_11_n_38 & n_1448));
 assign mul_109_11_n_242 = ~((n_79 | n_77) & (n_1177 | n_1183));
 assign mul_109_11_n_256 = ((n_1177 & ~n_81) | (n_79 & n_81));
 assign mul_109_11_n_255 = ((mul_109_11_n_39 & ~n_84) | (n_201 & n_84));
 assign n_224 = ~((n_83 | n_201) & (n_225 | mul_109_11_n_39));
 assign mul_109_11_n_245 = ~((n_82 & ~n_87) | (n_1195 & n_87));
 assign mul_109_11_n_247 = ~((n_88 & ~n_135) | (n_1176 & n_135));
 assign n_231 = ((n_229 & ~n_388) | (n_136 & n_388));
 assign mul_109_11_n_374 = ~((n_310 & ~n_1409) | (mul_109_11_n_19 & n_1409));
 assign mul_109_11_n_347 = ~((n_310 & ~n_1408) | (mul_109_11_n_19 & n_1408));
 assign mul_109_11_n_295 = ((mul_109_11_n_19 & ~n_1410) | (n_310 & n_1410));
 assign csa_tree_add_106_2_groupi_n_392 = ~((csa_tree_add_106_2_groupi_n_24 | n_203) & (n_213 | n_202));
 assign mul_109_11_n_303 = ~((n_31 | n_88) & (n_1196 | n_1176));
 assign mul_109_11_n_402 = ~(n_1449 & ~n_1382);
 assign csa_tree_add_106_2_groupi_n_411 = ~((csa_tree_add_106_2_groupi_n_9 | n_1178) & (csa_tree_add_106_2_groupi_n_17
    | n_1179));
 assign csa_tree_add_106_2_groupi_n_403 = ~((csa_tree_add_106_2_groupi_n_12 | n_1179) & (csa_tree_add_106_2_groupi_n_22
    | n_1178));
 assign csa_tree_add_106_2_groupi_n_399 = ~((csa_tree_add_106_2_groupi_n_64 | n_1179) & (csa_tree_add_106_2_groupi_n_51
    | n_1178));
 assign csa_tree_add_106_2_groupi_n_398 = ~((csa_tree_add_106_2_groupi_n_64 | n_1178) & (csa_tree_add_106_2_groupi_n_22
    | n_1179));
 assign csa_tree_add_106_2_groupi_n_397 = ~((csa_tree_add_106_2_groupi_n_65 | n_1178) & (csa_tree_add_106_2_groupi_n_62
    | n_1179));
 assign csa_tree_add_106_2_groupi_n_395 = ~((csa_tree_add_106_2_groupi_n_49 | n_1179) & (csa_tree_add_106_2_groupi_n_53
    | n_1178));
 assign csa_tree_add_106_2_groupi_n_394 = ~((csa_tree_add_106_2_groupi_n_62 | n_1178) & (csa_tree_add_106_2_groupi_n_51
    | n_1179));
 assign csa_tree_add_106_2_groupi_n_386 = ~((csa_tree_add_106_2_groupi_n_12 | n_1178) & (csa_tree_add_106_2_groupi_n_9
    | n_1179));
 assign csa_tree_add_106_2_groupi_n_353 = ~((csa_tree_add_106_2_groupi_n_65 | n_1179) & (csa_tree_add_106_2_groupi_n_49
    | n_1178));
 assign csa_tree_add_106_2_groupi_n_415 = ~((csa_tree_add_106_2_groupi_n_20 | n_203) & (csa_tree_add_106_2_groupi_n_24
    | n_202));
 assign csa_tree_add_106_2_groupi_n_417 = ~((n_365 | n_202) & (n_203 | n_209));
 assign csa_tree_add_106_2_groupi_n_391 = ~((csa_tree_add_106_2_groupi_n_31 | n_202) & (csa_tree_add_106_2_groupi_n_58
    | n_203));
 assign csa_tree_add_106_2_groupi_n_420 = ~((csa_tree_add_106_2_groupi_n_31 | n_203) & (csa_tree_add_106_2_groupi_n_52
    | n_202));
 assign csa_tree_add_106_2_groupi_n_404 = ~((n_202 | n_363) & (n_365 | n_203));
 assign csa_tree_add_106_2_groupi_n_423 = ~((csa_tree_add_106_2_groupi_n_19 | n_203) & (csa_tree_add_106_2_groupi_n_58
    | n_202));
 assign csa_tree_add_106_2_groupi_n_413 = ~((csa_tree_add_106_2_groupi_n_20 | n_202) & (csa_tree_add_106_2_groupi_n_52
    | n_203));
 assign n_259 = ((n_1326 | n_428) & (csa_tree_add_106_2_groupi_n_71 | n_322));
 assign n_232 = ~((n_136 & ~n_1409) | (n_229 & n_1409));
 assign mul_109_11_n_366 = ~((n_29 | n_88) & (n_1194 | n_1176));
 assign mul_109_11_n_367 = ~((n_26 | n_88) & (n_1193 | n_1176));
 assign mul_109_11_n_371 = ~((n_26 | n_310) & (n_1193 | mul_109_11_n_19));
 assign mul_109_11_n_370 = ~((n_29 | n_310) & (n_1194 | mul_109_11_n_19));
 assign mul_109_11_n_223 = ~((n_1452 | n_362) & (mul_109_11_n_52 | mul_109_11_n_38));
 assign mul_109_11_n_237 = ~((n_1454 | n_362) & (mul_109_11_n_31 | mul_109_11_n_38));
 assign mul_109_11_n_239 = ~((mul_109_11_n_41 & ~n_37) | (n_1143 & n_37));
 assign mul_109_11_n_140 = ~((n_1454 | n_106) & (mul_109_11_n_31 | n_749));
 assign mul_109_11_n_282 = ~((n_1450 | n_106) & (mul_109_11_n_56 | n_749));
 assign mul_109_11_n_207 = ~((n_1452 | n_106) & (mul_109_11_n_52 | n_749));
 assign mul_109_11_n_192 = ~((n_1452 | n_1) & (mul_109_11_n_52 | n_751));
 assign mul_109_11_n_275 = ~((n_1450 | n_1) & (mul_109_11_n_56 | n_751));
 assign mul_109_11_n_132 = ~((n_1454 | n_1) & (mul_109_11_n_31 | n_751));
 assign mul_109_11_n_250 = ~((mul_109_11_n_56 | n_433) & (n_1450 | n_777));
 assign mul_109_11_n_191 = ~((n_1452 | n_433) & (mul_109_11_n_52 | n_777));
 assign mul_109_11_n_133 = ~((n_1454 | n_433) & (mul_109_11_n_31 | n_777));
 assign mul_109_11_n_122 = ~((n_1454 | n_90) & (mul_109_11_n_31 | n_743));
 assign mul_109_11_n_177 = ~((n_1452 | n_90) & (mul_109_11_n_52 | n_743));
 assign mul_109_11_n_81 = ~((mul_109_11_n_52 | n_92) & (n_1452 | n_744));
 assign mul_109_11_n_121 = ~((n_1454 | n_92) & (mul_109_11_n_31 | n_744));
 assign mul_109_11_n_353 = ~((n_23 | n_88) & (n_1191 | n_1176));
 assign mul_109_11_n_352 = ~((n_24 | n_88) & (n_1192 | n_1176));
 assign mul_109_11_n_74 = ~((n_1454 | n_96) & (mul_109_11_n_31 | n_746));
 assign mul_109_11_n_109 = ~((n_1454 | n_95) & (mul_109_11_n_31 | n_745));
 assign mul_109_11_n_356 = ~((n_23 | n_310) & (n_1191 | mul_109_11_n_19));
 assign mul_109_11_n_357 = ~((n_24 | n_310) & (n_1192 | mul_109_11_n_19));
 assign n_234 = ~((n_1336 & n_403) | (n_1324 & n_404));
 assign n_1063 = ~((csa_tree_add_106_2_groupi_n_16 & n_393) | (n_1414 & n_395));
 assign n_1102 = ~((csa_tree_add_106_2_groupi_n_62 & n_160) | (n_1424 & n_402));
 assign n_1110 = ~((csa_tree_add_106_2_groupi_n_17 & n_416) | (n_1418 & n_418));
 assign n_1112 = ~((csa_tree_add_106_2_groupi_n_11 & n_416) | (n_1417 & n_418));
 assign n_1046 = ~((csa_tree_add_106_2_groupi_n_16 & n_160) | (n_1414 & n_402));
 assign n_1119 = ~((csa_tree_add_106_2_groupi_n_14 & n_416) | (n_1415 & n_418));
 assign n_1109 = ~((csa_tree_add_106_2_groupi_n_9 & n_416) | (n_1419 & n_418));
 assign n_1108 = ~((csa_tree_add_106_2_groupi_n_12 & n_416) | (n_1420 & n_418));
 assign n_1111 = ~((csa_tree_add_106_2_groupi_n_22 & n_416) | (n_1421 & n_418));
 assign n_1036 = ~((csa_tree_add_106_2_groupi_n_23 & n_421) | (n_1329 & n_422));
 assign n_1117 = ~((csa_tree_add_106_2_groupi_n_51 & n_416) | (n_1423 & n_418));
 assign n_1115 = ~((csa_tree_add_106_2_groupi_n_62 & n_416) | (n_1424 & n_418));
 assign n_1114 = ~((csa_tree_add_106_2_groupi_n_65 & n_416) | (n_1425 & n_418));
 assign n_1068 = ~((csa_tree_add_106_2_groupi_n_71 & n_421) | (n_1326 & n_422));
 assign n_1130 = ~((n_1331 & n_439) | (csa_tree_add_106_2_groupi_n_58 & n_104));
 assign n_1129 = ~((n_1332 & n_439) | (csa_tree_add_106_2_groupi_n_31 & n_104));
 assign n_1122 = ~((csa_tree_add_106_2_groupi_n_32 & n_104) | (n_1328 & n_439));
 assign n_1125 = ~((csa_tree_add_106_2_groupi_n_23 & n_104) | (n_1329 & n_439));
 assign n_1127 = ~((n_1335 & n_439) | (csa_tree_add_106_2_groupi_n_24 & n_104));
 assign n_1133 = ~((csa_tree_add_106_2_groupi_n_71 & n_104) | (n_1326 & n_439));
 assign n_1123 = ~((csa_tree_add_106_2_groupi_n_70 & n_104) | (n_1327 & n_439));
 assign n_1131 = ~((n_1330 & n_439) | (csa_tree_add_106_2_groupi_n_19 & n_104));
 assign n_1057 = ~((n_1335 & n_422) | (csa_tree_add_106_2_groupi_n_24 & n_421));
 assign n_1126 = ~((n_1334 & n_439) | (csa_tree_add_106_2_groupi_n_20 & n_104));
 assign n_1056 = ~((n_1334 & n_422) | (csa_tree_add_106_2_groupi_n_20 & n_421));
 assign n_1128 = ~((n_1333 & n_439) | (csa_tree_add_106_2_groupi_n_52 & n_104));
 assign n_1039 = ~((n_1330 & n_422) | (csa_tree_add_106_2_groupi_n_19 & n_421));
 assign n_1134 = ~((n_1335 & n_428) | (csa_tree_add_106_2_groupi_n_24 & n_322));
 assign n_1038 = ~((n_1331 & n_422) | (csa_tree_add_106_2_groupi_n_58 & n_421));
 assign n_1138 = ~((n_1334 & n_428) | (csa_tree_add_106_2_groupi_n_20 & n_322));
 assign n_1140 = ~((n_1330 & n_428) | (csa_tree_add_106_2_groupi_n_19 & n_322));
 assign n_1135 = ~((n_1331 & n_428) | (csa_tree_add_106_2_groupi_n_58 & n_322));
 assign n_1136 = ~((n_1332 & n_428) | (csa_tree_add_106_2_groupi_n_31 & n_322));
 assign n_1037 = ~((csa_tree_add_106_2_groupi_n_32 & n_421) | (n_1328 & n_422));
 assign n_1137 = ~((n_1333 & n_428) | (csa_tree_add_106_2_groupi_n_52 & n_322));
 assign n_1081 = ~((csa_tree_add_106_2_groupi_n_32 & n_322) | (n_1328 & n_428));
 assign n_925 = ~(n_129 | n_1170);
 assign n_1139 = ~((csa_tree_add_106_2_groupi_n_23 & n_322) | (n_1329 & n_428));
 assign n_1124 = ~((csa_tree_add_106_2_groupi_n_70 & n_322) | (n_1327 & n_428));
 assign n_1049 = ~((n_1332 & n_422) | (csa_tree_add_106_2_groupi_n_31 & n_421));
 assign n_924 = ~((n_428 & n_358) | (n_322 & n_209));
 assign n_1048 = ~((n_1333 & n_422) | (csa_tree_add_106_2_groupi_n_52 & n_421));
 assign n_830 = ~((n_67 & n_419) | (n_417 & n_1338));
 assign n_1035 = ~((csa_tree_add_106_2_groupi_n_70 & n_421) | (n_1327 & n_422));
 assign n_1066 = ~((n_402 & n_317) | (n_318 & n_160));
 assign n_876 = ~((n_358 & n_404) | (n_403 & n_209));
 assign n_1079 = ~(n_1325 ^ n_403);
 assign n_1067 = ~(n_1325 ^ n_421);
 assign n_1132 = ~(n_1325 ^ n_104);
 assign n_1113 = ~((csa_tree_add_106_2_groupi_n_13 & n_416) | (n_1416 & n_418));
 assign n_1059 = ~((csa_tree_add_106_2_groupi_n_69 & n_382) | (n_1412 & n_384));
 assign n_1033 = ~((csa_tree_add_106_2_groupi_n_68 & n_382) | (n_1413 & n_384));
 assign n_1074 = ~((n_1335 & n_404) | (csa_tree_add_106_2_groupi_n_24 & n_403));
 assign n_1044 = ~((csa_tree_add_106_2_groupi_n_14 & n_393) | (n_1415 & n_395));
 assign n_838 = ~((n_396 & n_67) | (n_394 & n_1338));
 assign csa_tree_mul_77_11_groupi_n_560 = ~(n_130 & (n_129 | n_137));
 assign n_889 = ~((n_364 | n_393) & (n_1180 | n_395));
 assign n_1344 = ~(csa_tree_mul_77_11_groupi_n_441 ^ csa_tree_mul_77_11_groupi_n_447);
 assign n_1096 = ~((csa_tree_add_106_2_groupi_n_13 & n_393) | (n_1416 & n_395));
 assign n_887 = ~((n_117 | n_382) & (n_214 | n_384));
 assign n_885 = ~((n_149 | n_382) & (n_1181 | n_384));
 assign n_1089 = ~((csa_tree_add_106_2_groupi_n_22 & n_382) | (n_1421 & n_384));
 assign n_1028 = ~((csa_tree_add_106_2_groupi_n_13 & n_160) | (n_1416 & n_402));
 assign n_1025 = ~((csa_tree_add_106_2_groupi_n_72 & n_160) | (n_1411 & n_402));
 assign n_1101 = ~((csa_tree_add_106_2_groupi_n_65 & n_160) | (n_1425 & n_402));
 assign n_886 = ~((n_119 | n_382) & (n_215 | n_384));
 assign n_750 = ~((n_136 & ~n_1410) | (n_229 & n_1410));
 assign n_1166 = ~(csa_tree_add_92_2_groupi_n_282 ^ n_6);
 assign n_1075 = ~((n_1330 & n_404) | (csa_tree_add_106_2_groupi_n_19 & n_403));
 assign n_1072 = ~((n_1331 & n_404) | (csa_tree_add_106_2_groupi_n_58 & n_403));
 assign n_1070 = ~((n_1333 & n_404) | (csa_tree_add_106_2_groupi_n_52 & n_403));
 assign n_843 = ~((n_439 & n_358) | (n_104 & n_209));
 assign n_1076 = ~((csa_tree_add_106_2_groupi_n_70 & n_403) | (n_1327 & n_404));
 assign n_719 = ~((n_31 | n_136) & (n_1196 | n_229));
 assign n_883 = ~((n_1337 | n_403) & (n_327 | n_404));
 assign n_1071 = ~((n_1332 & n_404) | (csa_tree_add_106_2_groupi_n_31 & n_403));
 assign n_1077 = ~((csa_tree_add_106_2_groupi_n_23 & n_403) | (n_1329 & n_404));
 assign n_1078 = ~((csa_tree_add_106_2_groupi_n_32 & n_403) | (n_1328 & n_404));
 assign n_1098 = ~((csa_tree_add_106_2_groupi_n_62 & n_393) | (n_1424 & n_395));
 assign n_1116 = ~((csa_tree_add_106_2_groupi_n_64 & n_416) | (n_1422 & n_418));
 assign n_1042 = ~((csa_tree_add_106_2_groupi_n_72 & n_416) | (n_1411 & n_418));
 assign n_1339 = ~(csa_tree_mul_77_11_groupi_n_582 ^ csa_tree_mul_77_11_groupi_n_507);
 assign n_882 = ~((n_377 | n_403) & (n_205 | n_404));
 assign n_1085 = ~((csa_tree_add_106_2_groupi_n_51 & n_382) | (n_1423 & n_384));
 assign n_880 = ~((n_355 | n_403) & (n_204 | n_404));
 assign n_1118 = ~((csa_tree_add_106_2_groupi_n_16 & n_416) | (n_1414 & n_418));
 assign n_1047 = ~((csa_tree_add_106_2_groupi_n_68 & n_160) | (n_1413 & n_402));
 assign n_1084 = ~((csa_tree_add_106_2_groupi_n_62 & n_382) | (n_1424 & n_384));
 assign n_881 = ~((n_350 | n_403) & (n_212 | n_404));
 assign n_1031 = ~((csa_tree_add_106_2_groupi_n_11 & n_160) | (n_1417 & n_402));
 assign n_1086 = ~((csa_tree_add_106_2_groupi_n_12 & n_382) | (n_1420 & n_384));
 assign n_872 = ~((n_375 | n_403) & (n_207 | n_404));
 assign n_1082 = ~((csa_tree_add_106_2_groupi_n_17 & n_382) | (n_1418 & n_384));
 assign n_845 = ~((n_382 | n_407) & (n_384 | n_1182));
 assign n_1061 = ~((csa_tree_add_106_2_groupi_n_11 & n_382) | (n_1417 & n_384));
 assign n_884 = ~((n_382 | n_364) & (n_384 | n_1180));
 assign n_888 = ~((n_407 | n_393) & (n_1182 | n_395));
 assign n_1120 = ~((csa_tree_add_106_2_groupi_n_13 & n_382) | (n_1416 & n_384));
 assign n_1087 = ~((csa_tree_add_106_2_groupi_n_9 & n_382) | (n_1419 & n_384));
 assign mul_109_11_n_364 = ~((n_26 | n_82) & (n_1193 | n_1195));
 assign n_1121 = ~((csa_tree_add_106_2_groupi_n_14 & n_382) | (n_1415 & n_384));
 assign n_1083 = ~((csa_tree_add_106_2_groupi_n_65 & n_382) | (n_1425 & n_384));
 assign n_759 = ~((n_29 | n_136) & (n_1194 | n_229));
 assign n_765 = ~((n_26 | n_136) & (n_1193 | n_229));
 assign n_1080 = ~((csa_tree_add_106_2_groupi_n_71 & n_403) | (n_1326 & n_404));
 assign n_1040 = ~((csa_tree_add_106_2_groupi_n_16 & n_382) | (n_1414 & n_384));
 assign n_1088 = ~((csa_tree_add_106_2_groupi_n_64 & n_382) | (n_1422 & n_384));
 assign n_1090 = ~((csa_tree_add_106_2_groupi_n_22 & n_393) | (n_1421 & n_395));
 assign n_1093 = ~((csa_tree_add_106_2_groupi_n_64 & n_393) | (n_1422 & n_395));
 assign n_1092 = ~((csa_tree_add_106_2_groupi_n_9 & n_393) | (n_1419 & n_395));
 assign n_1091 = ~((csa_tree_add_106_2_groupi_n_12 & n_393) | (n_1420 & n_395));
 assign n_1029 = ~((csa_tree_add_106_2_groupi_n_14 & n_160) | (n_1415 & n_402));
 assign n_1094 = ~((csa_tree_add_106_2_groupi_n_17 & n_393) | (n_1418 & n_395));
 assign n_1099 = ~((csa_tree_add_106_2_groupi_n_51 & n_393) | (n_1423 & n_395));
 assign n_1095 = ~((csa_tree_add_106_2_groupi_n_11 & n_393) | (n_1417 & n_395));
 assign n_1100 = ~((csa_tree_add_106_2_groupi_n_22 & n_160) | (n_1421 & n_402));
 assign n_1024 = ~((csa_tree_add_106_2_groupi_n_69 & n_160) | (n_1412 & n_402));
 assign n_1103 = ~((csa_tree_add_106_2_groupi_n_12 & n_160) | (n_1420 & n_402));
 assign n_728 = ~((n_23 | n_201) & (n_1191 | mul_109_11_n_39));
 assign n_1104 = ~((csa_tree_add_106_2_groupi_n_64 & n_160) | (n_1422 & n_402));
 assign n_841 = ~((n_385 & n_67) | (n_383 & n_1338));
 assign n_1105 = ~((csa_tree_add_106_2_groupi_n_51 & n_160) | (n_1423 & n_402));
 assign n_1064 = ~((csa_tree_add_106_2_groupi_n_68 & n_393) | (n_1413 & n_395));
 assign n_854 = ~((n_23 | n_82) & (n_1191 | n_1195));
 assign n_815 = ~((n_24 | n_82) & (n_1192 | n_1195));
 assign n_1060 = ~((csa_tree_add_106_2_groupi_n_72 & n_382) | (n_1411 & n_384));
 assign n_1106 = ~((csa_tree_add_106_2_groupi_n_9 & n_160) | (n_1419 & n_402));
 assign n_1097 = ~((csa_tree_add_106_2_groupi_n_65 & n_393) | (n_1425 & n_395));
 assign n_1052 = ~((csa_tree_add_106_2_groupi_n_69 & n_393) | (n_1412 & n_395));
 assign n_769 = ~((n_23 | n_136) & (n_1191 | n_229));
 assign n_770 = ~((n_24 | n_136) & (n_1192 | n_229));
 assign n_1107 = ~((csa_tree_add_106_2_groupi_n_17 & n_160) | (n_1418 & n_402));
 assign n_1053 = ~((csa_tree_add_106_2_groupi_n_72 & n_393) | (n_1411 & n_395));
 assign n_1073 = ~((n_1334 & n_404) | (csa_tree_add_106_2_groupi_n_20 & n_403));
 assign n_849 = ~((n_357 | n_104) & (n_439 | n_210));
 assign n_906 = ~((n_350 | n_104) & (n_212 | n_439));
 assign n_901 = ~((n_416 | n_149) & (n_418 | n_1181));
 assign n_809 = ~((n_416 | n_364) & (n_418 | n_1180));
 assign n_811 = ~((n_416 | n_407) & (n_418 | n_1182));
 assign n_898 = ~((n_364 | n_160) & (n_1180 | n_402));
 assign n_893 = ~((n_407 | n_160) & (n_1182 | n_402));
 assign n_899 = ~((n_149 | n_160) & (n_1181 | n_402));
 assign n_896 = ~((n_119 | n_160) & (n_215 | n_402));
 assign n_900 = ~((n_119 | n_416) & (n_215 | n_418));
 assign n_902 = ~((n_416 | n_117) & (n_418 | n_214));
 assign n_897 = ~((n_117 | n_160) & (n_214 | n_402));
 assign n_907 = ~((n_355 | n_104) & (n_204 | n_439));
 assign n_908 = ~((n_1337 | n_104) & (n_327 | n_439));
 assign n_909 = ~((n_377 | n_104) & (n_205 | n_439));
 assign n_910 = ~((n_375 | n_104) & (n_207 | n_439));
 assign n_850 = ~((n_349 | n_104) & (n_439 | n_211));
 assign n_241 = ~((csa_tree_add_106_2_groupi_n_11 | n_1178) & (csa_tree_add_106_2_groupi_n_13 | n_1179));
 assign n_240 = ~((csa_tree_add_106_2_groupi_n_16 | n_1179) & (csa_tree_add_106_2_groupi_n_14 | n_1178));
 assign n_239 = ~((csa_tree_add_106_2_groupi_n_16 | n_1178) & (csa_tree_add_106_2_groupi_n_68 | n_1179));
 assign n_238 = ~((csa_tree_add_106_2_groupi_n_11 | n_1179) & (csa_tree_add_106_2_groupi_n_17 | n_1178));
 assign n_237 = ~((csa_tree_add_106_2_groupi_n_13 | n_1178) & (csa_tree_add_106_2_groupi_n_14 | n_1179));
 assign n_1341 = ~(csa_tree_mul_77_11_groupi_n_566 ^ csa_tree_mul_77_11_groupi_n_571);
 assign n_236 = ~((n_202 | n_367) & (n_363 | n_203));
 assign n_1346 = ~(csa_tree_mul_77_11_groupi_n_367 ^ csa_tree_mul_77_11_groupi_n_406);
 assign n_1444 = ~(add_100_2_n_28 ^ add_100_2_n_19);
 assign n_1440 = ~(add_100_2_n_40 ^ add_100_2_n_17);
 assign n_1442 = ~(add_100_2_n_35 ^ add_100_2_n_13);
 assign n_1153 = ~(csa_tree_mul_77_11_groupi_n_617 ^ n_342);
 assign n_1340 = ~csa_tree_add_86_2_n_6;
 assign mul_109_11_n_85 = ~((n_100 | n_77) & (n_1197 | n_1183));
 assign n_1384 = ~(csa_tree_mul_77_11_groupi_n_592 ^ csa_tree_mul_77_11_groupi_n_508);
 assign n_235 = ~((mul_109_11_n_38 & n_201) | (n_362 & mul_109_11_n_39));
 assign n_230 = ~((mul_109_11_n_38 & n_82) | (n_362 & n_1195));
 assign n_228 = ~((mul_109_11_n_38 & n_136) | (n_362 & n_229));
 assign csa_tree_add_106_2_groupi_n_416 = ~((n_202 | n_152) & (n_203 | n_206));
 assign csa_tree_add_106_2_groupi_n_390 = ~((n_202 | n_206) & (n_213 | n_203));
 assign csa_tree_add_106_2_groupi_n_414 = ~((n_202 | n_208) & (n_203 | n_152));
 assign mul_109_11_n_234 = ~((mul_109_11_n_25 | n_74) & (n_1146 | n_1207));
 assign mul_109_11_n_224 = ~((n_60 | n_1184) & (n_1175 | n_11));
 assign csa_tree_add_106_2_groupi_n_412 = ~((n_207 | n_202) & (n_203 | n_208));
 assign mul_109_11_n_84 = ~((n_362 | n_77) & (mul_109_11_n_38 | n_1183));
 assign mul_109_11_n_190 = ~((n_1 | n_310) & (n_751 | mul_109_11_n_19));
 assign mul_109_11_n_189 = ~((n_433 | n_310) & (n_777 | mul_109_11_n_19));
 assign mul_109_11_n_159 = ~((n_106 | n_88) & (n_749 | n_1176));
 assign mul_109_11_n_173 = ~((n_433 | n_88) & (n_777 | n_1176));
 assign mul_109_11_n_174 = ~((n_1 | n_88) & (n_751 | n_1176));
 assign mul_109_11_n_208 = ~((n_310 | n_90) & (mul_109_11_n_19 | n_743));
 assign mul_109_11_n_209 = ~((n_310 | n_92) & (mul_109_11_n_19 | n_744));
 assign mul_109_11_n_135 = ~((n_106 | n_81) & (n_749 | n_1185));
 assign mul_109_11_n_193 = ~((n_90 | n_88) & (n_743 | n_1176));
 assign mul_109_11_n_194 = ~((n_92 | n_88) & (n_744 | n_1176));
 assign mul_109_11_n_108 = ~((n_310 | n_95) & (mul_109_11_n_19 | n_745));
 assign mul_109_11_n_102 = ~((n_310 | n_96) & (mul_109_11_n_19 | n_746));
 assign mul_109_11_n_335 = ~((n_19 | n_81) & (n_1189 | n_1185));
 assign mul_109_11_n_228 = ~((n_20 | n_81) & (n_1190 | n_1185));
 assign mul_109_11_n_123 = ~((n_106 | n_77) & (n_749 | n_1183));
 assign mul_109_11_n_147 = ~((n_1 | n_81) & (n_751 | n_1185));
 assign mul_109_11_n_146 = ~((n_433 | n_81) & (n_777 | n_1185));
 assign mul_109_11_n_214 = ~((n_95 | n_88) & (n_745 | n_1176));
 assign mul_109_11_n_215 = ~((n_96 | n_88) & (n_746 | n_1176));
 assign mul_109_11_n_340 = ~((n_19 | n_88) & (n_1189 | n_1176));
 assign mul_109_11_n_341 = ~((n_20 | n_88) & (n_1190 | n_1176));
 assign mul_109_11_n_137 = ~((n_1 | n_77) & (n_751 | n_1183));
 assign mul_109_11_n_136 = ~((n_433 | n_77) & (n_777 | n_1183));
 assign mul_109_11_n_119 = ~((n_106 | n_60) & (n_749 | n_1175));
 assign mul_109_11_n_361 = ~((n_310 | n_97) & (mul_109_11_n_19 | n_747));
 assign mul_109_11_n_161 = ~((n_310 | n_98) & (mul_109_11_n_19 | n_748));
 assign mul_109_11_n_162 = ~((n_90 | n_81) & (n_743 | n_1185));
 assign mul_109_11_n_163 = ~((n_92 | n_81) & (n_744 | n_1185));
 assign mul_109_11_n_345 = ~((n_19 | n_310) & (n_1189 | mul_109_11_n_19));
 assign mul_109_11_n_344 = ~((n_20 | n_310) & (n_1190 | mul_109_11_n_19));
 assign mul_109_11_n_105 = ~((n_106 | n_1146) & (n_749 | mul_109_11_n_25));
 assign mul_109_11_n_127 = ~((n_433 | n_60) & (n_777 | n_1175));
 assign mul_109_11_n_126 = ~((n_1 | n_60) & (n_751 | n_1175));
 assign mul_109_11_n_154 = ~((n_92 | n_77) & (n_744 | n_1183));
 assign mul_109_11_n_153 = ~((n_90 | n_77) & (n_743 | n_1183));
 assign mul_109_11_n_120 = ~((n_98 | n_88) & (n_748 | n_1176));
 assign mul_109_11_n_226 = ~((n_13 | n_77) & (n_1187 | n_1183));
 assign mul_109_11_n_318 = ~((n_12 | n_77) & (n_1186 | n_1183));
 assign mul_109_11_n_321 = ~((n_12 | n_81) & (n_1186 | n_1185));
 assign mul_109_11_n_320 = ~((n_13 | n_81) & (n_1187 | n_1185));
 assign mul_109_11_n_134 = ~((n_97 | n_88) & (n_747 | n_1176));
 assign mul_109_11_n_187 = ~((n_96 | n_81) & (n_746 | n_1185));
 assign mul_109_11_n_188 = ~((n_95 | n_81) & (n_745 | n_1185));
 assign mul_109_11_n_267 = ~((n_310 | n_99) & (mul_109_11_n_19 | n_1198));
 assign mul_109_11_n_296 = ~((n_60 | n_14) & (n_1175 | n_1188));
 assign mul_109_11_n_327 = ~((n_12 | n_88) & (n_1186 | n_1176));
 assign mul_109_11_n_328 = ~((n_13 | n_88) & (n_1187 | n_1176));
 assign mul_109_11_n_233 = ~((n_1194 | n_82) & (n_29 | n_1195));
 assign mul_109_11_n_268 = ~((n_310 | n_100) & (mul_109_11_n_19 | n_1197));
 assign mul_109_11_n_117 = ~((n_433 | n_1146) & (n_777 | mul_109_11_n_25));
 assign mul_109_11_n_301 = ~((n_11 | n_77) & (n_1184 | n_1183));
 assign mul_109_11_n_302 = ~((n_14 | n_77) & (n_1188 | n_1183));
 assign mul_109_11_n_332 = ~((n_310 | n_13) & (mul_109_11_n_19 | n_1187));
 assign mul_109_11_n_333 = ~((n_310 | n_12) & (mul_109_11_n_19 | n_1186));
 assign mul_109_11_n_372 = ~((n_1146 | n_73) & (mul_109_11_n_25 | n_1202));
 assign mul_109_11_n_307 = ~((n_11 | n_81) & (n_1184 | n_1185));
 assign mul_109_11_n_306 = ~((n_14 | n_81) & (n_1188 | n_1185));
 assign mul_109_11_n_83 = ~((n_1143 | n_75) & (mul_109_11_n_41 | n_1201));
 assign mul_109_11_n_206 = ~((n_1143 | n_101) & (mul_109_11_n_41 | n_1200));
 assign mul_109_11_n_272 = ~((n_60 | n_74) & (n_1175 | n_1207));
 assign mul_109_11_n_271 = ~((n_60 | n_73) & (n_1175 | n_1202));
 assign mul_109_11_n_118 = ~((n_1 | n_1146) & (n_751 | mul_109_11_n_25));
 assign mul_109_11_n_139 = ~((n_60 | n_92) & (n_1175 | n_744));
 assign mul_109_11_n_138 = ~((n_60 | n_90) & (n_1175 | n_743));
 assign mul_109_11_n_171 = ~((n_95 | n_77) & (n_745 | n_1183));
 assign mul_109_11_n_312 = ~((n_11 | n_88) & (n_1184 | n_1176));
 assign mul_109_11_n_313 = ~((n_14 | n_88) & (n_1188 | n_1176));
 assign mul_109_11_n_278 = ~((n_73 | n_77) & (n_1202 | n_1183));
 assign mul_109_11_n_279 = ~((n_74 | n_77) & (n_1207 | n_1183));
 assign mul_109_11_n_87 = ~((n_1146 | n_101) & (mul_109_11_n_25 | n_1200));
 assign mul_109_11_n_86 = ~((n_1146 | n_75) & (mul_109_11_n_25 | n_1201));
 assign mul_109_11_n_172 = ~((n_96 | n_77) & (n_746 | n_1183));
 assign mul_109_11_n_96 = ~((n_106 | n_1143) & (n_749 | mul_109_11_n_41));
 assign mul_109_11_n_168 = ~((n_1143 | n_100) & (mul_109_11_n_41 | n_1197));
 assign mul_109_11_n_167 = ~((n_1143 | n_99) & (mul_109_11_n_41 | n_1198));
 assign mul_109_11_n_317 = ~((n_310 | n_11) & (mul_109_11_n_19 | n_1184));
 assign mul_109_11_n_316 = ~((n_310 | n_14) & (mul_109_11_n_19 | n_1188));
 assign mul_109_11_n_285 = ~((n_74 | n_81) & (n_1207 | n_1185));
 assign mul_109_11_n_286 = ~((n_73 | n_81) & (n_1202 | n_1185));
 assign mul_109_11_n_151 = ~((n_60 | n_101) & (n_1175 | n_1200));
 assign mul_109_11_n_149 = ~((n_60 | n_75) & (n_1175 | n_1201));
 assign mul_109_11_n_277 = ~((n_99 | n_88) & (n_1198 | n_1176));
 assign mul_109_11_n_375 = ~((n_100 | n_88) & (n_1197 | n_1176));
 assign mul_109_11_n_196 = ~((n_1146 | n_100) & (mul_109_11_n_25 | n_1197));
 assign mul_109_11_n_195 = ~((n_1146 | n_99) & (mul_109_11_n_25 | n_1198));
 assign mul_109_11_n_322 = ~((n_75 | n_77) & (n_1201 | n_1183));
 assign mul_109_11_n_334 = ~((n_101 | n_77) & (n_1200 | n_1183));
 assign mul_109_11_n_210 = ~((n_97 | n_81) & (n_747 | n_1185));
 assign mul_109_11_n_211 = ~((n_98 | n_81) & (n_748 | n_1185));
 assign mul_109_11_n_144 = ~((n_1143 | n_98) & (mul_109_11_n_41 | n_748));
 assign mul_109_11_n_145 = ~((n_1143 | n_97) & (mul_109_11_n_41 | n_747));
 assign mul_109_11_n_298 = ~((n_73 | n_88) & (n_1202 | n_1176));
 assign mul_109_11_n_297 = ~((n_74 | n_88) & (n_1207 | n_1176));
 assign csa_tree_add_106_2_groupi_n_409 = ~((n_1178 | n_1181) & (n_1179 | n_214));
 assign csa_tree_add_106_2_groupi_n_405 = ~((n_1178 | n_1182) & (n_1179 | n_1180));
 assign csa_tree_add_106_2_groupi_n_402 = ~((n_1178 | n_1180) & (n_1179 | n_1181));
 assign csa_tree_add_106_2_groupi_n_389 = ~((n_1178 | n_214) & (n_215 | n_1179));
 assign csa_tree_add_106_2_groupi_n_418 = ~((n_327 | n_202) & (n_205 | n_203));
 assign csa_tree_add_106_2_groupi_n_393 = ~((n_202 | n_211) & (n_212 | n_203));
 assign csa_tree_add_106_2_groupi_n_425 = ~((n_212 | n_202) & (n_204 | n_203));
 assign csa_tree_add_106_2_groupi_n_401 = ~((n_202 | n_210) & (n_203 | n_211));
 assign csa_tree_add_106_2_groupi_n_424 = ~((n_204 | n_202) & (n_327 | n_203));
 assign csa_tree_add_106_2_groupi_n_421 = ~((n_205 | n_202) & (n_207 | n_203));
 assign mul_109_11_n_212 = ~((n_60 | n_99) & (n_1175 | n_1198));
 assign mul_109_11_n_213 = ~((n_60 | n_100) & (n_1175 | n_1197));
 assign mul_109_11_n_360 = ~((n_101 | n_81) & (n_1200 | n_1185));
 assign mul_109_11_n_346 = ~((n_75 | n_81) & (n_1201 | n_1185));
 assign mul_109_11_n_128 = ~((n_1146 | n_92) & (mul_109_11_n_25 | n_744));
 assign mul_109_11_n_129 = ~((n_1146 | n_90) & (mul_109_11_n_25 | n_743));
 assign mul_109_11_n_305 = ~((n_310 | n_73) & (mul_109_11_n_19 | n_1202));
 assign mul_109_11_n_304 = ~((n_310 | n_74) & (mul_109_11_n_19 | n_1207));
 assign mul_109_11_n_131 = ~((n_1143 | n_95) & (mul_109_11_n_41 | n_745));
 assign mul_109_11_n_130 = ~((n_1143 | n_96) & (mul_109_11_n_41 | n_746));
 assign mul_109_11_n_165 = ~((n_1146 | n_98) & (mul_109_11_n_25 | n_748));
 assign mul_109_11_n_164 = ~((n_1146 | n_97) & (mul_109_11_n_25 | n_747));
 assign mul_109_11_n_221 = ~((n_99 | n_77) & (n_1198 | n_1183));
 assign mul_109_11_n_157 = ~((n_60 | n_96) & (n_1175 | n_746));
 assign mul_109_11_n_158 = ~((n_60 | n_95) & (n_1175 | n_745));
 assign mul_109_11_n_103 = ~((n_1143 | n_433) & (mul_109_11_n_41 | n_777));
 assign n_227 = ~((n_24 & mul_109_11_n_39) | (n_1192 & n_201));
 assign mul_109_11_n_104 = ~((n_1 | n_1143) & (n_751 | mul_109_11_n_41));
 assign mul_109_11_n_287 = ~((n_310 | n_75) & (mul_109_11_n_19 | n_1201));
 assign mul_109_11_n_184 = ~((n_60 | n_97) & (n_1175 | n_747));
 assign mul_109_11_n_183 = ~((n_60 | n_98) & (n_1175 | n_748));
 assign mul_109_11_n_281 = ~((n_101 | n_88) & (n_1200 | n_1176));
 assign mul_109_11_n_280 = ~((n_75 | n_88) & (n_1201 | n_1176));
 assign mul_109_11_n_115 = ~((n_1143 | n_92) & (mul_109_11_n_41 | n_744));
 assign mul_109_11_n_116 = ~((n_1143 | n_90) & (mul_109_11_n_41 | n_743));
 assign mul_109_11_n_112 = ~((n_100 | n_81) & (n_1197 | n_1185));
 assign mul_109_11_n_110 = ~((n_99 | n_81) & (n_1198 | n_1185));
 assign mul_109_11_n_143 = ~((n_1146 | n_96) & (mul_109_11_n_25 | n_746));
 assign mul_109_11_n_142 = ~((n_1146 | n_95) & (mul_109_11_n_25 | n_745));
 assign mul_109_11_n_288 = ~((n_310 | n_101) & (mul_109_11_n_19 | n_1200));
 assign mul_109_11_n_200 = ~((n_98 | n_77) & (n_748 | n_1183));
 assign mul_109_11_n_199 = ~((n_97 | n_77) & (n_747 | n_1183));
 assign n_867 = ~((n_19 | n_82) & (n_1189 | n_1195));
 assign n_754 = ~((n_75 | n_136) & (n_1201 | n_229));
 assign n_869 = ~((n_75 | n_82) & (n_1201 | n_1195));
 assign n_868 = ~((n_101 | n_82) & (n_1200 | n_1195));
 assign n_735 = ~((n_100 | n_201) & (n_1197 | mul_109_11_n_39));
 assign n_738 = ~((n_99 | n_201) & (n_1198 | mul_109_11_n_39));
 assign n_736 = ~((n_101 | n_201) & (n_1200 | mul_109_11_n_39));
 assign n_721 = ~((n_75 | n_201) & (n_1201 | mul_109_11_n_39));
 assign n_859 = ~((n_99 | n_82) & (n_1198 | n_1195));
 assign n_858 = ~((n_100 | n_82) & (n_1197 | n_1195));
 assign n_891 = ~((n_119 | n_393) & (n_215 | n_395));
 assign n_775 = ~((n_74 | n_136) & (n_1207 | n_229));
 assign n_755 = ~((n_73 | n_136) & (n_1202 | n_229));
 assign n_860 = ~((n_74 | n_82) & (n_1207 | n_1195));
 assign n_861 = ~((n_73 | n_82) & (n_1202 | n_1195));
 assign n_729 = ~((n_74 | n_201) & (n_1207 | mul_109_11_n_39));
 assign n_722 = ~((n_73 | n_201) & (n_1202 | mul_109_11_n_39));
 assign n_762 = ~((n_11 | n_136) & (n_1184 | n_229));
 assign n_776 = ~((n_14 | n_136) & (n_1188 | n_229));
 assign n_857 = ~((n_14 | n_82) & (n_1188 | n_1195));
 assign n_865 = ~((n_11 | n_82) & (n_1184 | n_1195));
 assign n_760 = ~((n_99 | n_136) & (n_1198 | n_229));
 assign n_761 = ~((n_100 | n_136) & (n_1197 | n_229));
 assign n_730 = ~((n_14 | n_201) & (n_1188 | mul_109_11_n_39));
 assign n_725 = ~((n_11 | n_201) & (n_1184 | mul_109_11_n_39));
 assign n_771 = ~((n_13 | n_136) & (n_1187 | n_229));
 assign n_756 = ~((n_12 | n_136) & (n_1186 | n_229));
 assign n_737 = ~((n_98 | n_201) & (n_748 | mul_109_11_n_39));
 assign n_742 = ~((n_97 | n_201) & (n_747 | mul_109_11_n_39));
 assign n_856 = ~((n_13 | n_82) & (n_1187 | n_1195));
 assign n_864 = ~((n_12 | n_82) & (n_1186 | n_1195));
 assign n_870 = ~((n_98 | n_82) & (n_748 | n_1195));
 assign n_871 = ~((n_97 | n_82) & (n_747 | n_1195));
 assign n_726 = ~((n_12 | n_201) & (n_1186 | mul_109_11_n_39));
 assign n_723 = ~((n_13 | n_201) & (n_1187 | mul_109_11_n_39));
 assign n_817 = ~((n_153 | n_421) & (n_206 | n_422));
 assign n_818 = ~((n_421 | n_242) & (n_422 | n_152));
 assign n_825 = ~((n_154 | n_421) & (n_213 | n_422));
 assign n_903 = ~((n_154 | n_104) & (n_213 | n_439));
 assign n_904 = ~((n_153 | n_104) & (n_206 | n_439));
 assign n_753 = ~((n_98 | n_136) & (n_748 | n_229));
 assign n_764 = ~((n_97 | n_136) & (n_747 | n_229));
 assign n_741 = ~((n_96 | n_201) & (n_746 | mul_109_11_n_39));
 assign n_731 = ~((n_95 | n_201) & (n_745 | mul_109_11_n_39));
 assign n_905 = ~((n_242 | n_104) & (n_152 | n_439));
 assign n_772 = ~((n_19 | n_136) & (n_1189 | n_229));
 assign n_757 = ~((n_20 | n_136) & (n_1190 | n_229));
 assign n_879 = ~((n_154 | n_403) & (n_213 | n_404));
 assign n_877 = ~((n_153 | n_403) & (n_206 | n_404));
 assign n_862 = ~((n_95 | n_82) & (n_745 | n_1195));
 assign n_863 = ~((n_96 | n_82) & (n_746 | n_1195));
 assign n_874 = ~((n_242 | n_403) & (n_152 | n_404));
 assign n_819 = ~((n_421 | n_170) & (n_422 | n_208));
 assign n_911 = ~((n_170 | n_104) & (n_208 | n_439));
 assign n_758 = ~((n_101 | n_136) & (n_1200 | n_229));
 assign n_866 = ~((n_20 | n_82) & (n_1190 | n_1195));
 assign n_724 = ~((n_19 | n_201) & (n_1189 | mul_109_11_n_39));
 assign n_740 = ~((n_92 | n_201) & (n_744 | mul_109_11_n_39));
 assign n_739 = ~((n_90 | n_201) & (n_743 | mul_109_11_n_39));
 assign n_727 = ~((n_20 | n_201) & (n_1190 | mul_109_11_n_39));
 assign n_767 = ~((n_95 | n_136) & (n_745 | n_229));
 assign n_763 = ~((n_96 | n_136) & (n_746 | n_229));
 assign n_895 = ~((n_90 | n_82) & (n_743 | n_1195));
 assign n_855 = ~((n_92 | n_82) & (n_744 | n_1195));
 assign n_873 = ~((n_170 | n_403) & (n_208 | n_404));
 assign n_921 = ~((n_154 | n_322) & (n_213 | n_428));
 assign n_916 = ~((n_153 | n_322) & (n_206 | n_428));
 assign n_915 = ~((n_322 | n_242) & (n_428 | n_152));
 assign n_820 = ~((n_1337 | n_421) & (n_327 | n_422));
 assign n_732 = ~((n_433 | n_201) & (n_777 | mul_109_11_n_39));
 assign n_734 = ~((n_1 | n_201) & (n_751 | mul_109_11_n_39));
 assign n_853 = ~((n_1 | n_82) & (n_751 | n_1195));
 assign n_894 = ~((n_433 | n_82) & (n_777 | n_1195));
 assign n_766 = ~((n_92 | n_136) & (n_744 | n_229));
 assign n_768 = ~((n_90 | n_136) & (n_743 | n_229));
 assign n_821 = ~((n_1324 | n_1471) & (n_1336 | n_243));
 assign n_822 = ~((n_377 | n_421) & (n_205 | n_422));
 assign n_823 = ~((n_375 | n_421) & (n_207 | n_422));
 assign n_923 = ~((n_357 | n_322) & (n_428 | n_210));
 assign n_733 = ~((n_106 | n_201) & (n_749 | mul_109_11_n_39));
 assign n_804 = ~((n_106 | n_82) & (n_749 | n_1195));
 assign n_773 = ~((n_1 | n_136) & (n_751 | n_229));
 assign n_774 = ~((n_433 | n_136) & (n_777 | n_229));
 assign n_824 = ~((n_355 | n_421) & (n_204 | n_422));
 assign n_922 = ~((n_322 | n_349) & (n_428 | n_211));
 assign n_919 = ~((n_1337 | n_322) & (n_327 | n_428));
 assign n_752 = ~((n_106 | n_136) & (n_749 | n_229));
 assign n_832 = ~((n_350 | n_421) & (n_212 | n_422));
 assign n_917 = ~((n_355 | n_322) & (n_204 | n_428));
 assign n_920 = ~((n_350 | n_322) & (n_212 | n_428));
 assign n_222 = ~((csa_tree_add_92_2_groupi_n_207 & ~n_1370) | (n_223 & n_1370));
 assign n_837 = ~((n_394 | n_69) & (n_396 | n_244));
 assign n_840 = ~((n_69 | n_383) & (n_244 | n_385));
 assign n_828 = ~((n_69 | n_417) & (n_244 | n_419));
 assign n_914 = ~((n_170 | n_322) & (n_208 | n_428));
 assign mul_109_11_n_169 = ~((n_749 | n_310) & (n_106 | mul_109_11_n_19));
 assign n_918 = ~((n_377 | n_322) & (n_205 | n_428));
 assign n_913 = ~((n_375 | n_322) & (n_207 | n_428));
 assign n_834 = ~((n_421 | n_357) & (n_422 | n_210));
 assign n_835 = ~((n_421 | n_349) & (n_422 | n_211));
 assign n_875 = ~((n_357 | n_403) & (n_210 | n_404));
 assign n_878 = ~((n_349 | n_403) & (n_211 | n_404));
 assign n_892 = ~((n_117 | n_393) & (n_214 | n_395));
 assign n_890 = ~((n_149 | n_393) & (n_1181 | n_395));
 assign csa_tree_add_92_2_groupi_n_65 = (n_4 ^ n_3);
 assign csa_tree_add_86_2_n_6 = ~(csa_tree_mul_77_11_groupi_n_567 ^ csa_tree_mul_77_11_groupi_n_581);
 assign n_1069 = ~(n_443 ^ n_120);
 assign n_1016 = ~(n_1401 ^ n_1371);
 assign csa_tree_add_106_2_groupi_n_45 = ~({in1[0]} ^ {in2[0]});
 assign n_1381 = ~n_1382;
 assign n_1459 = ~(csa_tree_mul_77_11_groupi_n_453 & csa_tree_mul_77_11_groupi_n_475);
 assign csa_tree_add_86_2_n_165 = ~(csa_tree_add_86_2_n_17 | n_8);
 assign csa_tree_add_86_2_n_146 = ~(csa_tree_add_86_2_n_30 | n_8);
 assign csa_tree_add_86_2_n_155 = ~(csa_tree_add_86_2_n_14 | n_8);
 assign csa_tree_add_86_2_n_45 = ~(csa_tree_add_86_2_n_19 | n_431);
 assign csa_tree_mul_77_11_groupi_n_498 = ~(n_325 & n_166);
 assign csa_tree_mul_77_11_groupi_n_495 = ~(n_251 & n_250);
 assign csa_tree_add_86_2_n_379 = ~(csa_tree_add_86_2_n_34 | n_401);
 assign csa_tree_add_86_2_n_114 = ~(csa_tree_add_86_2_n_15 | n_114);
 assign csa_tree_add_86_2_n_320 = ~(n_1336 | ~n_2);
 assign csa_tree_add_86_2_n_208 = ~(csa_tree_add_86_2_n_10 | n_114);
 assign n_1460 = ~(n_83 & n_82);
 assign csa_tree_add_86_2_n_55 = ~(csa_tree_add_86_2_n_19 | n_8);
 assign csa_tree_add_86_2_n_202 = ~(csa_tree_add_86_2_n_9 | n_114);
 assign n_277 = ~(csa_tree_mul_77_11_groupi_n_476 & csa_tree_mul_77_11_groupi_n_525);
 assign csa_tree_add_86_2_n_205 = ~(csa_tree_add_86_2_n_19 | n_114);
 assign n_1461 = ~(n_374 & stall);
 assign csa_tree_add_86_2_n_378 = ~(csa_tree_add_86_2_n_23 | n_401);
 assign csa_tree_add_86_2_n_138 = ~(csa_tree_add_86_2_n_8 | n_431);
 assign n_1462 = (n_3 | n_4);
 assign csa_tree_add_86_2_n_89 = ~(csa_tree_add_86_2_n_8 | n_8);
 assign n_1463 = ~(csa_tree_mul_77_11_groupi_n_526 | csa_tree_mul_77_11_groupi_n_504);
 assign csa_tree_mul_77_11_groupi_n_419 = (n_339 & n_340);
 assign csa_tree_add_86_2_n_116 = ~(csa_tree_add_86_2_n_16 | n_8);
 assign csa_tree_add_86_2_n_376 = ~(n_401 | n_405);
 assign csa_tree_add_86_2_n_48 = ~(csa_tree_add_86_2_n_10 | n_8);
 assign csa_tree_add_86_2_n_368 = ~(csa_tree_add_86_2_n_8 | n_401);
 assign mul_109_11_n_329 = ~(n_310 & ~{out1[0]});
 assign csa_tree_add_86_2_n_197 = ~(csa_tree_add_86_2_n_30 | n_114);
 assign csa_tree_add_86_2_n_102 = ~(csa_tree_add_86_2_n_16 | n_431);
 assign csa_tree_add_86_2_n_46 = ~(csa_tree_add_86_2_n_9 | n_431);
 assign csa_tree_add_86_2_n_39 = ~(csa_tree_add_86_2_n_15 | n_431);
 assign csa_tree_add_86_2_n_99 = ~(csa_tree_add_86_2_n_17 | n_431);
 assign csa_tree_add_86_2_n_194 = ~(csa_tree_add_86_2_n_15 | n_376);
 assign csa_tree_add_86_2_n_142 = ~(csa_tree_add_86_2_n_19 | n_420);
 assign csa_tree_add_86_2_n_118 = ~(csa_tree_add_86_2_n_30 | n_426);
 assign csa_tree_add_86_2_n_183 = ~(csa_tree_add_86_2_n_9 | n_426);
 assign csa_tree_mul_77_11_groupi_n_428 = ~(n_341 | ~n_339);
 assign csa_tree_add_86_2_n_78 = ~(csa_tree_add_86_2_n_23 | n_376);
 assign csa_tree_mul_77_11_groupi_n_386 = ~(n_252 | n_341);
 assign csa_tree_add_86_2_n_185 = ~(csa_tree_add_86_2_n_9 | n_409);
 assign csa_tree_add_86_2_n_247 = ~(n_401 | n_351);
 assign csa_tree_add_86_2_n_120 = ~(csa_tree_add_86_2_n_14 | n_409);
 assign csa_tree_add_86_2_n_97 = ~(csa_tree_add_86_2_n_15 | n_409);
 assign csa_tree_add_86_2_n_201 = ~(csa_tree_add_86_2_n_9 | n_376);
 assign csa_tree_mul_77_11_groupi_n_554 = ~(n_130 & ~n_129);
 assign csa_tree_add_86_2_n_277 = ~(n_1336 | ~n_113);
 assign mul_109_11_n_384 = (n_370 | mul_109_11_n_19);
 assign csa_tree_add_86_2_n_200 = ~(csa_tree_add_86_2_n_16 | n_420);
 assign csa_tree_mul_77_11_groupi_n_448 = ~(n_343 & ~n_438);
 assign n_1464 = ~(csa_tree_mul_77_11_groupi_n_476 | csa_tree_mul_77_11_groupi_n_525);
 assign csa_tree_add_86_2_n_136 = ~(csa_tree_add_86_2_n_30 | n_376);
 assign csa_tree_add_86_2_n_190 = ~(n_405 | n_376);
 assign csa_tree_add_86_2_n_159 = ~(csa_tree_add_86_2_n_19 | n_376);
 assign csa_tree_add_86_2_n_145 = ~(csa_tree_add_86_2_n_17 | n_376);
 assign csa_tree_add_86_2_n_130 = ~(csa_tree_add_86_2_n_8 | n_376);
 assign csa_tree_add_86_2_n_49 = ~(csa_tree_add_86_2_n_8 | n_409);
 assign csa_tree_add_86_2_n_211 = ~(csa_tree_add_86_2_n_17 | n_114);
 assign csa_tree_add_86_2_n_203 = ~(csa_tree_add_86_2_n_16 | n_114);
 assign csa_tree_add_86_2_n_168 = ~(csa_tree_add_86_2_n_8 | n_114);
 assign csa_tree_add_86_2_n_177 = ~(csa_tree_add_86_2_n_14 | n_114);
 assign csa_tree_add_86_2_n_53 = ~(csa_tree_add_86_2_n_17 | n_409);
 assign csa_tree_add_86_2_n_242 = ~(csa_tree_add_86_2_n_19 | n_401);
 assign csa_tree_add_86_2_n_152 = ~(csa_tree_add_86_2_n_10 | n_376);
 assign csa_tree_add_86_2_n_213 = ~(n_420 | n_405);
 assign csa_tree_add_86_2_n_170 = ~(csa_tree_add_86_2_n_34 | n_409);
 assign csa_tree_add_86_2_n_63 = ~(csa_tree_add_86_2_n_16 | n_409);
 assign csa_tree_add_86_2_n_93 = ~(csa_tree_add_86_2_n_16 | n_426);
 assign csa_tree_add_86_2_n_176 = ~(csa_tree_add_86_2_n_34 | n_376);
 assign csa_tree_add_86_2_n_87 = ~(csa_tree_add_86_2_n_14 | n_376);
 assign csa_tree_add_86_2_n_100 = ~(csa_tree_add_86_2_n_23 | n_114);
 assign csa_tree_add_86_2_n_377 = ~(csa_tree_add_86_2_n_17 | n_401);
 assign csa_tree_add_86_2_n_375 = ~(csa_tree_add_86_2_n_16 | n_401);
 assign csa_tree_add_86_2_n_370 = ~(csa_tree_add_86_2_n_10 | n_401);
 assign csa_tree_add_86_2_n_367 = ~(n_401 | n_434);
 assign csa_tree_add_86_2_n_366 = ~(csa_tree_add_86_2_n_9 | n_401);
 assign csa_tree_add_86_2_n_79 = ~(csa_tree_add_86_2_n_23 | n_409);
 assign csa_tree_add_86_2_n_363 = ~(csa_tree_add_86_2_n_15 | n_401);
 assign csa_tree_add_86_2_n_252 = ~(n_1336 | ~n_406);
 assign csa_tree_add_86_2_n_50 = ~(csa_tree_add_86_2_n_10 | n_409);
 assign csa_tree_add_86_2_n_167 = ~(csa_tree_add_86_2_n_19 | n_409);
 assign csa_tree_add_86_2_n_123 = ~(csa_tree_add_86_2_n_30 | n_409);
 assign csa_tree_add_86_2_n_206 = ~(csa_tree_add_86_2_n_16 | n_376);
 assign n_1155 = (n_1401 | n_1371);
 assign n_1206 = ~(n_61 & n_77);
 assign n_233 = ~(n_1413 & n_418);
 assign n_1149 = (n_443 | n_120);
 assign n_1382 = ~(n_1450 | n_362);
 assign n_219 = ~n_220;
 assign n_217 = ~n_218;
 assign csa_tree_add_86_2_n_180 = ~(csa_tree_add_86_2_n_34 | n_8);
 assign csa_tree_add_86_2_n_149 = ~(csa_tree_add_86_2_n_14 | n_431);
 assign csa_tree_add_86_2_n_160 = ~(csa_tree_add_86_2_n_23 | n_431);
 assign csa_tree_add_86_2_n_51 = ~(csa_tree_add_86_2_n_34 | n_114);
 assign n_1467 = ~(n_341 & stall);
 assign csa_tree_add_86_2_n_387 = ~(csa_tree_add_86_2_n_9 | n_420);
 assign csa_tree_add_86_2_n_384 = ~(csa_tree_add_86_2_n_34 | n_420);
 assign csa_tree_add_86_2_n_225 = ~(csa_tree_add_86_2_n_14 | n_420);
 assign csa_tree_add_86_2_n_221 = ~(csa_tree_add_86_2_n_17 | n_420);
 assign csa_tree_add_86_2_n_195 = ~(n_420 | n_434);
 assign csa_tree_add_86_2_n_181 = ~(csa_tree_add_86_2_n_10 | n_420);
 assign csa_tree_add_86_2_n_178 = ~(csa_tree_add_86_2_n_15 | n_420);
 assign csa_tree_add_86_2_n_143 = ~(csa_tree_add_86_2_n_23 | n_420);
 assign csa_tree_add_86_2_n_113 = ~(csa_tree_add_86_2_n_8 | n_420);
 assign mul_109_11_n_381 = ~(mul_109_11_n_38 | n_311);
 assign csa_tree_add_86_2_n_62 = ~(csa_tree_add_86_2_n_8 | n_426);
 assign csa_tree_add_86_2_n_65 = ~(csa_tree_add_86_2_n_10 | n_426);
 assign csa_tree_add_86_2_n_119 = ~(csa_tree_add_86_2_n_15 | n_426);
 assign csa_tree_add_86_2_n_193 = ~(csa_tree_add_86_2_n_19 | n_426);
 assign mul_109_11_n_403 = ~(mul_109_11_n_38 | n_800);
 assign csa_tree_add_86_2_n_271 = ~(n_1336 | ~n_425);
 assign csa_tree_add_86_2_n_196 = ~(csa_tree_add_86_2_n_14 | n_426);
 assign csa_tree_add_86_2_n_80 = ~(csa_tree_add_86_2_n_23 | n_426);
 assign csa_tree_add_86_2_n_117 = ~(csa_tree_add_86_2_n_17 | n_426);
 assign csa_tree_add_86_2_n_71 = ~(csa_tree_add_86_2_n_34 | n_426);
 assign mul_109_11_n_376 = ~(mul_109_11_n_38 | n_86);
 assign csa_tree_mul_77_11_groupi_n_509 = ~(n_374 | ~n_131);
 assign csa_tree_add_86_2_n_38 = ~(n_208 | n_376);
 assign csa_tree_add_86_2_n_92 = ~(csa_tree_add_86_2_n_23 | n_8);
 assign csa_tree_add_86_2_n_104 = ~(n_206 | n_426);
 assign csa_tree_add_86_2_n_298 = ~(n_1336 | ~n_430);
 assign csa_tree_add_86_2_n_187 = ~(csa_tree_add_86_2_n_34 | n_431);
 assign csa_tree_add_86_2_n_112 = ~(csa_tree_add_86_2_n_30 | n_431);
 assign csa_tree_add_86_2_n_212 = ~(n_114 | n_152);
 assign csa_tree_add_86_2_n_199 = ~(n_213 | n_420);
 assign csa_tree_add_86_2_n_69 = ~(n_206 | n_376);
 assign csa_tree_mul_77_11_groupi_n_553 = ~(n_148 | ~n_137);
 assign csa_tree_add_86_2_n_128 = ~(n_213 | n_376);
 assign csa_tree_add_86_2_n_121 = ~(n_213 | n_114);
 assign csa_tree_mul_77_11_groupi_n_510 = ~(n_151 & n_150);
 assign csa_tree_add_86_2_n_108 = ~(n_420 | n_208);
 assign csa_tree_add_86_2_n_90 = ~(n_114 | n_206);
 assign csa_tree_add_86_2_n_204 = ~(csa_tree_add_86_2_n_15 | n_8);
 assign csa_tree_add_86_2_n_386 = ~(n_420 | n_152);
 assign n_1466 = ~(csa_tree_mul_77_11_groupi_n_407 & csa_tree_mul_77_11_groupi_n_369);
 assign csa_tree_add_86_2_n_210 = ~(csa_tree_add_86_2_n_9 | n_8);
 assign csa_tree_add_86_2_n_96 = ~(csa_tree_add_86_2_n_10 | n_431);
 assign n_1465 = ~(csa_tree_mul_77_11_groupi_n_526 & csa_tree_mul_77_11_groupi_n_504);
 assign csa_tree_add_86_2_n_129 = ~(n_213 | n_426);
 assign csa_tree_add_86_2_n_115 = ~(n_213 | n_431);
 assign csa_tree_add_86_2_n_385 = ~(n_420 | n_206);
 assign csa_tree_add_86_2_n_163 = ~(n_213 | n_409);
 assign csa_tree_add_86_2_n_209 = ~(n_376 | n_152);
 assign csa_tree_add_86_2_n_380 = ~(n_401 | n_208);
 assign csa_tree_add_86_2_n_373 = ~(n_401 | n_206);
 assign csa_tree_add_86_2_n_361 = ~(n_401 | n_152);
 assign csa_tree_add_86_2_n_103 = ~(n_206 | n_8);
 assign csa_tree_add_86_2_n_137 = ~(n_213 | n_8);
 assign csa_tree_add_86_2_n_381 = ~(n_213 | n_401);
 assign n_220 = ~(n_229 & n_1468);
 assign n_1205 = ~(n_61 | n_77);
 assign n_1156 = ~(n_1401 & n_1371);
 assign n_1150 = ~(n_443 & n_120);
 assign n_1170 = ~(n_265 & ~n_148);
 assign n_1168 = ~(n_412 | n_1476);
 assign n_1034 = ~(n_362 | n_88);
 assign n_218 = ~(mul_109_11_n_38 | n_1176);
 assign n_1209 = ~(n_362 & n_81);
 assign n_1208 = ~(n_362 | n_81);
 assign n_1203 = ~(n_362 | n_60);
 assign n_1204 = ~(n_362 & n_60);
 assign n_1163 = ~(n_136 & n_135);
 assign csa_tree_mul_77_11_groupi_n_521 = ~(n_264 | n_374);
 assign n_276 = ~(n_114 | n_434);
 assign n_272 = ~(n_420 | n_351);
 assign n_270 = ~(n_405 | n_114);
 assign n_271 = ~(n_8 | n_152);
 assign n_263 = ~(n_409 | n_208);
 assign n_269 = ~(n_434 | n_426);
 assign n_275 = ~(n_405 | n_8);
 assign n_274 = ({in1[0]} & {in2[0]});
 assign n_1383 = ~(n_114 | n_208);
 assign n_1378 = ~(n_8 | n_208);
 assign n_273 = ~(n_431 | n_152);
 assign n_268 = ~(n_376 | n_434);
 assign n_260 = ~(n_208 | n_426);
 assign n_267 = ~(n_405 | n_426);
 assign n_266 = ~(n_409 | n_152);
 assign n_262 = ~(n_206 | n_431);
 assign n_261 = ~(n_409 | n_206);
 assign n_1430 = ~(n_426 | n_152);
 assign n_1158 = ~n_91;
 assign csa_tree_add_86_2_n_28 = ~{in5[6]};
 assign csa_tree_add_106_2_groupi_n_21 = ~n_1348;
 assign n_1157 = ~n_94;
 assign csa_tree_add_86_2_n_27 = ~{in5[5]};
 assign csa_tree_add_86_2_n_26 = ~{in5[1]};
 assign n_265 = ~csa_tree_mul_77_11_groupi_n_594;
 assign csa_tree_add_86_2_n_5 = ~{in5[0]};
 assign n_250 = ~n_325;
 assign n_791 = ~n_324;
 assign n_1473 = ~n_342;
 assign csa_tree_add_86_2_n_3 = ~{in5[4]};
 assign csa_tree_add_106_2_groupi_n_46 = ~n_1447;
 assign n_797 = ~n_347;
 assign n_264 = ~n_150;
 assign n_798 = ~n_321;
 assign mul_109_11_n_26 = ~n_370;
 assign n_1177 = ~n_79;
 assign n_209 = ~n_359;
 assign n_244 = ~n_69;
 assign n_1196 = ~n_31;
 assign n_1194 = ~n_29;
 assign n_1182 = ~n_407;
 assign n_211 = ~n_349;
 assign n_212 = ~n_350;
 assign n_1192 = ~n_24;
 assign n_205 = ~n_377;
 assign n_204 = ~n_355;
 assign n_215 = ~n_119;
 assign n_1180 = ~n_364;
 assign n_1337 = ~n_327;
 assign n_1189 = ~n_19;
 assign n_1190 = ~n_20;
 assign n_1188 = ~n_14;
 assign n_1184 = ~n_11;
 assign n_208 = ~n_170;
 assign n_206 = ~n_153;
 assign n_213 = ~n_154;
 assign n_242 = ~n_152;
 assign n_1207 = ~n_74;
 assign n_1200 = ~n_101;
 assign n_1201 = ~n_75;
 assign n_1178 = ~csa_tree_add_106_2_groupi_n_335;
 assign n_202 = ~csa_tree_add_106_2_groupi_n_337;
 assign n_203 = ~csa_tree_add_106_2_groupi_n_227;
 assign n_1179 = ~csa_tree_add_106_2_groupi_n_229;
 assign n_1471 = ~n_422;
 assign n_1478 = ~n_414;
 assign n_1470 = ~n_412;
 assign n_748 = ~n_98;
 assign n_1476 = ~n_416;
 assign n_747 = ~n_97;
 assign n_800 = ~mul_109_11_n_393;
 assign n_743 = ~n_90;
 assign n_749 = ~n_106;
 assign n_1143 = ~mul_109_11_n_41;
 assign n_1146 = ~mul_109_11_n_25;
 assign n_1175 = ~n_60;
 assign n_1183 = ~n_77;
 assign n_1195 = ~n_82;
 assign csa_tree_add_86_2_n_29 = ~{in5[7]};
 assign csa_tree_add_106_2_groupi_n_15 = ~n_1349;
 assign n_223 = ~csa_tree_add_92_2_groupi_n_207;
 assign n_252 = ~n_444;
 assign n_251 = ~n_166;
 assign csa_tree_add_86_2_n_4 = ~{in5[3]};
 assign csa_tree_add_86_2_n_25 = ~{in5[2]};
 assign n_1338 = ~n_76;
 assign n_1468 = ~n_135;
 assign n_709 = ~n_71;
 assign n_557 = ~n_15;
 assign n_225 = ~n_83;
 assign n_1199 = ~n_34;
 assign csa_tree_add_106_2_groupi_n_48 = ~n_1347;
 assign n_1477 = ~n_415;
 assign n_1193 = ~n_26;
 assign n_207 = ~n_375;
 assign n_1336 = ~n_1324;
 assign n_1191 = ~n_23;
 assign n_214 = ~n_117;
 assign n_1181 = ~n_149;
 assign n_210 = ~n_357;
 assign n_1186 = ~n_12;
 assign n_1187 = ~n_13;
 assign n_1202 = ~n_73;
 assign n_1198 = ~n_99;
 assign n_1197 = ~n_100;
 assign n_1474 = ~n_86;
 assign n_745 = ~n_95;
 assign n_746 = ~n_96;
 assign n_243 = ~n_421;
 assign n_744 = ~n_92;
 assign n_777 = ~n_433;
 assign n_751 = ~n_1;
 assign n_1472 = ~n_311;
 assign mul_109_11_n_38 = ~n_362;
 assign n_1185 = ~n_81;
 assign n_201 = ~mul_109_11_n_39;
 assign n_1176 = ~n_88;
 assign n_229 = ~n_136;
 assign mul_109_11_n_19 = ~n_310;
 assign n_465 = ~stall;
 assign mul_74_11_n_28 = ~(mul_74_11_n_27 & mul_74_11_n_464);
 assign n_1294 = ~(mul_74_11_n_570 ^ mul_74_11_n_462);
 assign mul_74_11_n_570 = ((mul_74_11_n_568 & mul_74_11_n_480) | ((mul_74_11_n_480 & mul_74_11_n_449)
    | (mul_74_11_n_449 & mul_74_11_n_568)));
 assign n_1295 = (mul_74_11_n_480 ^ (mul_74_11_n_449 ^ mul_74_11_n_568));
 assign mul_74_11_n_568 = ((mul_74_11_n_566 & mul_74_11_n_492) | ((mul_74_11_n_492 & mul_74_11_n_481)
    | (mul_74_11_n_481 & mul_74_11_n_566)));
 assign n_1296 = (mul_74_11_n_492 ^ (mul_74_11_n_481 ^ mul_74_11_n_566));
 assign mul_74_11_n_566 = ((mul_74_11_n_561 & mul_74_11_n_509) | ((mul_74_11_n_509 & mul_74_11_n_493)
    | (mul_74_11_n_493 & mul_74_11_n_561)));
 assign n_1297 = (mul_74_11_n_509 ^ (mul_74_11_n_493 ^ mul_74_11_n_561));
 assign n_1298 = (mul_74_11_n_564 ^ mul_74_11_n_524);
 assign mul_74_11_n_564 = ~(mul_74_11_n_538 & (mul_74_11_n_560 | mul_74_11_n_535));
 assign n_1299 = ~(mul_74_11_n_560 ^ mul_74_11_n_546);
 assign n_1300 = (mul_74_11_n_559 ^ mul_74_11_n_545);
 assign mul_74_11_n_561 = ~(mul_74_11_n_558 & (mul_74_11_n_548 | mul_74_11_n_552));
 assign mul_74_11_n_560 = ~(mul_74_11_n_551 | (mul_74_11_n_555 & mul_74_11_n_547));
 assign mul_74_11_n_559 = ~(mul_74_11_n_532 & (mul_74_11_n_554 | mul_74_11_n_537));
 assign mul_74_11_n_558 = ~(mul_74_11_n_542 | (mul_74_11_n_556 | (mul_74_11_n_551 & mul_74_11_n_549)));
 assign n_1301 = (mul_74_11_n_555 ^ mul_74_11_n_540);
 assign mul_74_11_n_556 = ~(mul_74_11_n_517 & (mul_74_11_n_550 | mul_74_11_n_552));
 assign mul_74_11_n_554 = ~mul_74_11_n_555;
 assign mul_74_11_n_555 = ~(mul_74_11_n_550 & mul_74_11_n_548);
 assign n_1302 = (mul_74_11_n_539 ^ mul_74_11_n_531);
 assign mul_74_11_n_552 = ~(mul_74_11_n_547 & mul_74_11_n_549);
 assign mul_74_11_n_551 = ~(mul_74_11_n_534 & (mul_74_11_n_532 | mul_74_11_n_533));
 assign mul_74_11_n_550 = ~(mul_74_11_n_543 | (mul_74_11_n_536 & mul_74_11_n_513));
 assign mul_74_11_n_549 = ~(mul_74_11_n_535 | mul_74_11_n_516);
 assign mul_74_11_n_548 = ~(mul_74_11_n_512 & mul_74_11_n_536);
 assign mul_74_11_n_547 = ~(mul_74_11_n_537 | mul_74_11_n_533);
 assign mul_74_11_n_546 = ~(mul_74_11_n_535 | ~mul_74_11_n_538);
 assign mul_74_11_n_545 = ~(mul_74_11_n_533 | ~mul_74_11_n_534);
 assign n_1303 = ~(mul_74_11_n_523 ^ mul_74_11_n_518);
 assign mul_74_11_n_543 = ~(mul_74_11_n_526 & (mul_74_11_n_525 | mul_74_11_n_506));
 assign mul_74_11_n_542 = ~(mul_74_11_n_538 | mul_74_11_n_516);
 assign n_1304 = (mul_74_11_n_522 ^ mul_74_11_n_503);
 assign mul_74_11_n_540 = ~(mul_74_11_n_537 | ~mul_74_11_n_532);
 assign mul_74_11_n_539 = ~(mul_74_11_n_506 & (mul_74_11_n_523 | mul_74_11_n_505));
 assign mul_74_11_n_538 = ~(mul_74_11_n_508 & mul_74_11_n_529);
 assign mul_74_11_n_537 = ~(mul_74_11_n_528 | mul_74_11_n_519);
 assign mul_74_11_n_536 = ~(mul_74_11_n_525 | mul_74_11_n_505);
 assign mul_74_11_n_535 = ~(mul_74_11_n_508 | mul_74_11_n_529);
 assign mul_74_11_n_534 = ~(mul_74_11_n_530 & mul_74_11_n_527);
 assign mul_74_11_n_533 = ~(mul_74_11_n_530 | mul_74_11_n_527);
 assign mul_74_11_n_532 = ~(mul_74_11_n_528 & mul_74_11_n_519);
 assign mul_74_11_n_531 = ~(mul_74_11_n_525 | ~mul_74_11_n_526);
 assign mul_74_11_n_529 = ((mul_74_11_n_461 & mul_74_11_n_470) | ((mul_74_11_n_470 & mul_74_11_n_394)
    | (mul_74_11_n_394 & mul_74_11_n_461)));
 assign mul_74_11_n_530 = (mul_74_11_n_470 ^ (mul_74_11_n_394 ^ mul_74_11_n_461));
 assign mul_74_11_n_527 = ((mul_74_11_n_478 & mul_74_11_n_471) | ((mul_74_11_n_471 & mul_74_11_n_392)
    | (mul_74_11_n_392 & mul_74_11_n_478)));
 assign mul_74_11_n_528 = (mul_74_11_n_471 ^ (mul_74_11_n_392 ^ mul_74_11_n_478));
 assign mul_74_11_n_526 = ~(mul_74_11_n_520 & mul_74_11_n_485);
 assign mul_74_11_n_525 = ~(mul_74_11_n_520 | mul_74_11_n_485);
 assign mul_74_11_n_524 = ~(mul_74_11_n_516 | ~mul_74_11_n_517);
 assign mul_74_11_n_523 = ~(mul_74_11_n_512 | mul_74_11_n_513);
 assign mul_74_11_n_522 = ~(mul_74_11_n_491 & (mul_74_11_n_502 | mul_74_11_n_490));
 assign mul_74_11_n_519 = ((mul_74_11_n_454 & mul_74_11_n_479) | ((mul_74_11_n_479 & mul_74_11_n_409)
    | (mul_74_11_n_409 & mul_74_11_n_454)));
 assign mul_74_11_n_520 = (mul_74_11_n_479 ^ (mul_74_11_n_409 ^ mul_74_11_n_454));
 assign mul_74_11_n_518 = ~(mul_74_11_n_505 | ~mul_74_11_n_506);
 assign mul_74_11_n_517 = ~(mul_74_11_n_510 & mul_74_11_n_507);
 assign mul_74_11_n_516 = ~(mul_74_11_n_510 | mul_74_11_n_507);
 assign mul_74_11_n_513 = ~(mul_74_11_n_500 & (mul_74_11_n_499 | mul_74_11_n_491));
 assign mul_74_11_n_512 = ~(mul_74_11_n_502 | mul_74_11_n_504);
 assign n_1306 = ~(mul_74_11_n_496 ^ mul_74_11_n_28);
 assign mul_74_11_n_509 = ((mul_74_11_n_468 & mul_74_11_n_420) | ((mul_74_11_n_420 & mul_74_11_n_446)
    | (mul_74_11_n_446 & mul_74_11_n_468)));
 assign mul_74_11_n_510 = (mul_74_11_n_420 ^ (mul_74_11_n_446 ^ mul_74_11_n_468));
 assign mul_74_11_n_507 = ((mul_74_11_n_460 & mul_74_11_n_469) | ((mul_74_11_n_469 & mul_74_11_n_407)
    | (mul_74_11_n_407 & mul_74_11_n_460)));
 assign mul_74_11_n_508 = (mul_74_11_n_469 ^ (mul_74_11_n_407 ^ mul_74_11_n_460));
 assign mul_74_11_n_506 = ~(mul_74_11_n_484 & mul_74_11_n_476);
 assign mul_74_11_n_505 = ~(mul_74_11_n_484 | mul_74_11_n_476);
 assign mul_74_11_n_504 = ~(mul_74_11_n_489 & (n_1503 | mul_74_11_n_465));
 assign mul_74_11_n_503 = ~(mul_74_11_n_499 | ~mul_74_11_n_500);
 assign mul_74_11_n_501 = ~mul_74_11_n_502;
 assign mul_74_11_n_502 = ~(mul_74_11_n_495 | mul_74_11_n_497);
 assign mul_74_11_n_500 = ~(n_1503 & mul_74_11_n_465);
 assign mul_74_11_n_499 = ~(n_1503 | mul_74_11_n_465);
 assign mul_74_11_n_498 = ~(mul_74_11_n_491 & ~mul_74_11_n_490);
 assign mul_74_11_n_497 = ~(mul_74_11_n_27 & (mul_74_11_n_25 | mul_74_11_n_26));
 assign mul_74_11_n_496 = ~(mul_74_11_n_450 & (mul_74_11_n_483 | mul_74_11_n_451));
 assign mul_74_11_n_495 = ~(mul_74_11_n_477 & (mul_74_11_n_25 | mul_74_11_n_456));
 assign mul_74_11_n_492 = ((mul_74_11_n_445 & mul_74_11_n_419) | ((mul_74_11_n_419 & mul_74_11_n_405)
    | (mul_74_11_n_405 & mul_74_11_n_445)));
 assign mul_74_11_n_493 = (mul_74_11_n_419 ^ (mul_74_11_n_405 ^ mul_74_11_n_445));
 assign mul_74_11_n_491 = ~(mul_74_11_n_23 & mul_74_11_n_441);
 assign mul_74_11_n_490 = ~mul_74_11_n_489;
 assign mul_74_11_n_489 = (mul_74_11_n_23 | mul_74_11_n_441);
 assign mul_74_11_n_485 = ~(mul_74_11_n_439 & (mul_74_11_n_24 | mul_74_11_n_443));
 assign mul_74_11_n_484 = (mul_74_11_n_24 ^ mul_74_11_n_455);
 assign mul_74_11_n_483 = ~mul_74_11_n_482;
 assign mul_74_11_n_480 = ((mul_74_11_n_404 & mul_74_11_n_413) | ((mul_74_11_n_413 & mul_74_11_n_226)
    | (mul_74_11_n_226 & mul_74_11_n_404)));
 assign mul_74_11_n_481 = (mul_74_11_n_413 ^ (mul_74_11_n_226 ^ mul_74_11_n_404));
 assign mul_74_11_n_478 = ((mul_74_11_n_386 & mul_74_11_n_16) | ((mul_74_11_n_16 & mul_74_11_n_400) |
    (mul_74_11_n_400 & mul_74_11_n_386)));
 assign mul_74_11_n_479 = (mul_74_11_n_16 ^ (mul_74_11_n_400 ^ mul_74_11_n_386));
 assign mul_74_11_n_477 = ~(mul_74_11_n_464 & ~mul_74_11_n_450);
 assign mul_74_11_n_482 = ~(mul_74_11_n_456 & mul_74_11_n_26);
 assign mul_74_11_n_476 = ~(mul_74_11_n_429 & (mul_74_11_n_438 | mul_74_11_n_434));
 assign mul_74_11_n_470 = ((mul_74_11_n_408 & mul_74_11_n_390) | ((mul_74_11_n_390 & mul_74_11_n_380)
    | (mul_74_11_n_380 & mul_74_11_n_408)));
 assign mul_74_11_n_471 = (mul_74_11_n_390 ^ (mul_74_11_n_380 ^ mul_74_11_n_408));
 assign mul_74_11_n_468 = ((mul_74_11_n_384 & mul_74_11_n_393) | ((mul_74_11_n_393 & mul_74_11_n_270)
    | (mul_74_11_n_270 & mul_74_11_n_384)));
 assign mul_74_11_n_469 = (mul_74_11_n_393 ^ (mul_74_11_n_270 ^ mul_74_11_n_384));
 assign mul_74_11_n_472 = ~(mul_74_11_n_458 & mul_74_11_n_414);
 assign n_1309 = (mul_74_11_n_34 ^ mul_74_11_n_453);
 assign mul_74_11_n_465 = ~(mul_74_11_n_457 & mul_74_11_n_21);
 assign mul_74_11_n_462 = ~(mul_74_11_n_448 ^ mul_74_11_n_374);
 assign mul_74_11_n_464 = ~(mul_74_11_n_440 & mul_74_11_n_417);
 assign mul_74_11_n_460 = ((mul_74_11_n_391 & mul_74_11_n_389) | ((mul_74_11_n_389 & mul_74_11_n_379)
    | (mul_74_11_n_379 & mul_74_11_n_391)));
 assign mul_74_11_n_461 = (mul_74_11_n_389 ^ (mul_74_11_n_379 ^ mul_74_11_n_391));
 assign mul_74_11_n_459 = ~(mul_74_11_n_450 & ~mul_74_11_n_451);
 assign mul_74_11_n_458 = ~(mul_74_11_n_453 & mul_74_11_n_403);
 assign mul_74_11_n_457 = ~(mul_74_11_n_422 & mul_74_11_n_418);
 assign mul_74_11_n_456 = ~(mul_74_11_n_444 | mul_74_11_n_431);
 assign mul_74_11_n_455 = ~((mul_74_11_n_424 & ~mul_74_11_n_436) | (mul_74_11_n_401 & mul_74_11_n_436));
 assign mul_74_11_n_454 = ~(mul_74_11_n_430 & (mul_74_11_n_435 | mul_74_11_n_382));
 assign mul_74_11_n_448 = ((mul_74_11_n_412 & mul_74_11_n_93) | ((mul_74_11_n_93 & mul_74_11_n_310) |
    (mul_74_11_n_310 & mul_74_11_n_412)));
 assign mul_74_11_n_449 = (mul_74_11_n_93 ^ (mul_74_11_n_310 ^ mul_74_11_n_412));
 assign mul_74_11_n_453 = ((mul_74_11_n_410 & mul_74_11_n_377) | ((mul_74_11_n_377 & mul_74_11_n_269)
    | (mul_74_11_n_269 & mul_74_11_n_410)));
 assign n_1310 = (mul_74_11_n_377 ^ (mul_74_11_n_269 ^ mul_74_11_n_410));
 assign mul_74_11_n_445 = ((mul_74_11_n_406 & mul_74_11_n_211) | ((mul_74_11_n_211 & mul_74_11_n_271)
    | (mul_74_11_n_271 & mul_74_11_n_406)));
 assign mul_74_11_n_446 = (mul_74_11_n_211 ^ (mul_74_11_n_271 ^ mul_74_11_n_406));
 assign mul_74_11_n_444 = ~(mul_74_11_n_432 | mul_74_11_n_414);
 assign mul_74_11_n_443 = ~(mul_74_11_n_436 | mul_74_11_n_424);
 assign mul_74_11_n_452 = ~(mul_74_11_n_433 & ~mul_74_11_n_431);
 assign mul_74_11_n_451 = ~(mul_74_11_n_416 | mul_74_11_n_425);
 assign mul_74_11_n_450 = ~(mul_74_11_n_416 & mul_74_11_n_425);
 assign mul_74_11_n_439 = ~(mul_74_11_n_436 & mul_74_11_n_424);
 assign mul_74_11_n_442 = (mul_74_11_n_15 ^ mul_74_11_n_421);
 assign mul_74_11_n_441 = ~((mul_74_11_n_398 & mul_74_11_n_17) | ((mul_74_11_n_17 & n_1505) | (n_1505
    & mul_74_11_n_398)));
 assign mul_74_11_n_440 = (mul_74_11_n_17 ^ mul_74_11_n_19);
 assign mul_74_11_n_438 = ~mul_74_11_n_437;
 assign mul_74_11_n_436 = ((mul_74_11_n_385 & mul_74_11_n_370) | ((mul_74_11_n_370 & mul_74_11_n_260)
    | (mul_74_11_n_260 & mul_74_11_n_385)));
 assign mul_74_11_n_437 = (mul_74_11_n_370 ^ (mul_74_11_n_260 ^ mul_74_11_n_385));
 assign mul_74_11_n_435 = ~(mul_74_11_n_402 | mul_74_11_n_372);
 assign mul_74_11_n_434 = ~(mul_74_11_n_423 | mul_74_11_n_421);
 assign mul_74_11_n_433 = ~mul_74_11_n_432;
 assign mul_74_11_n_432 = ~(mul_74_11_n_426 | mul_74_11_n_364);
 assign mul_74_11_n_431 = ~(mul_74_11_n_427 | mul_74_11_n_396);
 assign mul_74_11_n_430 = ~(mul_74_11_n_402 & mul_74_11_n_372);
 assign mul_74_11_n_429 = ~(mul_74_11_n_423 & mul_74_11_n_421);
 assign mul_74_11_n_428 = ~((mul_74_11_n_415 & ~mul_74_11_n_381) | (mul_74_11_n_395 & mul_74_11_n_381));
 assign mul_74_11_n_427 = ~mul_74_11_n_426;
 assign mul_74_11_n_424 = ~mul_74_11_n_401;
 assign mul_74_11_n_423 = ~mul_74_11_n_15;
 assign mul_74_11_n_425 = ((mul_74_11_n_14 & mul_74_11_n_262) | ((mul_74_11_n_262 & mul_74_11_n_315)
    | (mul_74_11_n_315 & mul_74_11_n_14)));
 assign mul_74_11_n_426 = (mul_74_11_n_262 ^ (mul_74_11_n_315 ^ mul_74_11_n_14));
 assign mul_74_11_n_419 = ((mul_74_11_n_264 & mul_74_11_n_290) | ((mul_74_11_n_290 & mul_74_11_n_345)
    | (mul_74_11_n_345 & mul_74_11_n_264)));
 assign mul_74_11_n_420 = (mul_74_11_n_290 ^ (mul_74_11_n_345 ^ mul_74_11_n_264));
 assign mul_74_11_n_421 = ((mul_74_11_n_10 & mul_74_11_n_343) | ((mul_74_11_n_343 & mul_74_11_n_261)
    | (mul_74_11_n_261 & mul_74_11_n_10)));
 assign mul_74_11_n_422 = (mul_74_11_n_343 ^ (mul_74_11_n_261 ^ mul_74_11_n_10));
 assign mul_74_11_n_418 = ~(mul_74_11_n_381 & mul_74_11_n_415);
 assign mul_74_11_n_417 = ~(mul_74_11_n_22 | mul_74_11_n_13);
 assign mul_74_11_n_416 = (mul_74_11_n_399 ^ mul_74_11_n_387);
 assign mul_74_11_n_415 = ~mul_74_11_n_395;
 assign mul_74_11_n_412 = ((mul_74_11_n_265 & mul_74_11_n_92) | ((mul_74_11_n_92 & mul_74_11_n_355) |
    (mul_74_11_n_355 & mul_74_11_n_265)));
 assign mul_74_11_n_413 = (mul_74_11_n_92 ^ (mul_74_11_n_355 ^ mul_74_11_n_265));
 assign mul_74_11_n_410 = ((mul_74_11_n_362 & mul_74_11_n_318) | ((mul_74_11_n_318 & mul_74_11_n_204)
    | (mul_74_11_n_204 & mul_74_11_n_362)));
 assign n_1311 = (mul_74_11_n_318 ^ (mul_74_11_n_204 ^ mul_74_11_n_362));
 assign mul_74_11_n_408 = ((mul_74_11_n_267 & mul_74_11_n_90) | ((mul_74_11_n_90 & mul_74_11_n_344) |
    (mul_74_11_n_344 & mul_74_11_n_267)));
 assign mul_74_11_n_409 = (mul_74_11_n_90 ^ (mul_74_11_n_344 ^ mul_74_11_n_267));
 assign mul_74_11_n_406 = ((mul_74_11_n_346 & mul_74_11_n_212) | ((mul_74_11_n_212 & mul_74_11_n_8) |
    (mul_74_11_n_8 & mul_74_11_n_346)));
 assign mul_74_11_n_407 = (mul_74_11_n_212 ^ (mul_74_11_n_8 ^ mul_74_11_n_346));
 assign mul_74_11_n_404 = ((mul_74_11_n_266 & mul_74_11_n_227) | ((mul_74_11_n_227 & mul_74_11_n_354)
    | (mul_74_11_n_354 & mul_74_11_n_266)));
 assign mul_74_11_n_405 = (mul_74_11_n_227 ^ (mul_74_11_n_354 ^ mul_74_11_n_266));
 assign mul_74_11_n_403 = (mul_74_11_n_383 | mul_74_11_n_378);
 assign mul_74_11_n_414 = ~(mul_74_11_n_383 & mul_74_11_n_378);
 assign mul_74_11_n_400 = ~(mul_74_11_n_369 & (mul_74_11_n_366 | mul_74_11_n_287));
 assign mul_74_11_n_402 = ~(mul_74_11_n_368 & (mul_74_11_n_367 | mul_74_11_n_285));
 assign mul_74_11_n_401 = ~(mul_74_11_n_11 ^ mul_74_11_n_286);
 assign mul_74_11_n_398 = ~mul_74_11_n_397;
 assign mul_74_11_n_396 = ~mul_74_11_n_364;
 assign mul_74_11_n_397 = ((mul_74_11_n_316 & mul_74_11_n_289) | ((mul_74_11_n_289 & mul_74_11_n_258)
    | (mul_74_11_n_258 & mul_74_11_n_316)));
 assign mul_74_11_n_399 = (mul_74_11_n_289 ^ (mul_74_11_n_258 ^ mul_74_11_n_316));
 assign mul_74_11_n_393 = ((mul_74_11_n_348 & mul_74_11_n_210) | ((mul_74_11_n_210 & mul_74_11_n_259)
    | (mul_74_11_n_259 & mul_74_11_n_348)));
 assign mul_74_11_n_394 = (mul_74_11_n_210 ^ (mul_74_11_n_259 ^ mul_74_11_n_348));
 assign mul_74_11_n_391 = ((mul_74_11_n_347 & mul_74_11_n_257) | ((mul_74_11_n_257 & mul_74_11_n_263)
    | (mul_74_11_n_263 & mul_74_11_n_347)));
 assign mul_74_11_n_392 = (mul_74_11_n_257 ^ (mul_74_11_n_263 ^ mul_74_11_n_347));
 assign mul_74_11_n_395 = ~(mul_74_11_n_388 & mul_74_11_n_357);
 assign mul_74_11_n_389 = ((mul_74_11_n_291 & n_1292) | ((n_1292 & mul_74_11_n_91) | (mul_74_11_n_91
    & mul_74_11_n_291)));
 assign mul_74_11_n_390 = (n_1292 ^ (mul_74_11_n_91 ^ mul_74_11_n_291));
 assign mul_74_11_n_388 = ~(mul_74_11_n_312 & (mul_74_11_n_324 | mul_74_11_n_323));
 assign mul_74_11_n_387 = ~((mul_74_11_n_371 & ~mul_74_11_n_280) | (mul_74_11_n_342 & mul_74_11_n_280));
 assign mul_74_11_n_386 = ~(mul_74_11_n_375 & mul_74_11_n_339);
 assign mul_74_11_n_385 = ~(mul_74_11_n_335 & (mul_74_11_n_334 | mul_74_11_n_325));
 assign mul_74_11_n_384 = ~((mul_74_11_n_282 | mul_74_11_n_340) & (mul_74_11_n_311 | n_1292));
 assign mul_74_11_n_383 = ~((mul_74_11_n_275 & ~n_1504) | (mul_74_11_n_276 & n_1504));
 assign mul_74_11_n_382 = ~((mul_74_11_n_327 & ~mul_74_11_n_9) | (mul_74_11_n_328 & mul_74_11_n_9));
 assign mul_74_11_n_380 = ~(mul_74_11_n_331 & (mul_74_11_n_332 | mul_74_11_n_288));
 assign mul_74_11_n_379 = ~(mul_74_11_n_281 ^ mul_74_11_n_349);
 assign mul_74_11_n_381 = (mul_74_11_n_12 ^ mul_74_11_n_325);
 assign mul_74_11_n_378 = (mul_74_11_n_317 & mul_74_11_n_231);
 assign mul_74_11_n_377 = (mul_74_11_n_317 ^ mul_74_11_n_231);
 assign mul_74_11_n_376 = ~(mul_74_11_n_280 | ~mul_74_11_n_371);
 assign mul_74_11_n_375 = ~(mul_74_11_n_328 & (mul_74_11_n_273 | mul_74_11_n_84));
 assign mul_74_11_n_374 = ~(mul_74_11_n_350 ^ mul_74_11_n_310);
 assign mul_74_11_n_373 = ~((mul_74_11_n_321 & ~mul_74_11_n_351) | (mul_74_11_n_322 & mul_74_11_n_351));
 assign mul_74_11_n_371 = ~mul_74_11_n_342;
 assign mul_74_11_n_372 = (mul_74_11_n_268 & mul_74_11_n_230);
 assign mul_74_11_n_370 = (mul_74_11_n_268 ^ mul_74_11_n_230);
 assign mul_74_11_n_369 = ~(mul_74_11_n_274 & mul_74_11_n_353);
 assign mul_74_11_n_368 = ~(mul_74_11_n_352 & mul_74_11_n_322);
 assign mul_74_11_n_367 = ~(mul_74_11_n_352 | mul_74_11_n_322);
 assign mul_74_11_n_366 = ~(mul_74_11_n_274 | mul_74_11_n_353);
 assign n_1312 = ~(mul_74_11_n_362 | (mul_74_11_n_329 & mul_74_11_n_184));
 assign mul_74_11_n_364 = ~(mul_74_11_n_360 & mul_74_11_n_336);
 assign mul_74_11_n_360 = ~(mul_74_11_n_333 & ~mul_74_11_n_326);
 assign mul_74_11_n_357 = ~(mul_74_11_n_324 & mul_74_11_n_323);
 assign mul_74_11_n_356 = ~((mul_74_11_n_35 & ~mul_74_11_n_277) | (n_1292 & mul_74_11_n_277));
 assign mul_74_11_n_355 = ~(mul_74_11_n_314 | (mul_74_11_n_6 & n_1286));
 assign mul_74_11_n_362 = ~(mul_74_11_n_329 | mul_74_11_n_184);
 assign mul_74_11_n_354 = ~(mul_74_11_n_313 & ~(mul_74_11_n_6 & mul_74_11_n_138));
 assign mul_74_11_n_352 = ~mul_74_11_n_351;
 assign mul_74_11_n_350 = ~(mul_74_11_n_292 ^ mul_74_11_n_94);
 assign mul_74_11_n_349 = ~((n_1292 & ~mul_74_11_n_311) | (mul_74_11_n_35 & mul_74_11_n_311));
 assign mul_74_11_n_348 = ~((mul_74_11_n_309 | mul_74_11_n_156) & (mul_74_11_n_240 | mul_74_11_n_143));
 assign mul_74_11_n_347 = ~(mul_74_11_n_341 & ~(mul_74_11_n_239 & mul_74_11_n_155));
 assign mul_74_11_n_346 = ~((mul_74_11_n_309 | mul_74_11_n_143) & (mul_74_11_n_240 | mul_74_11_n_153));
 assign mul_74_11_n_353 = ~(mul_74_11_n_4 & mul_74_11_n_296);
 assign mul_74_11_n_345 = ~(mul_74_11_n_295 & ~(mul_74_11_n_6 & mul_74_11_n_154));
 assign mul_74_11_n_344 = ~(mul_74_11_n_320 & mul_74_11_n_308);
 assign mul_74_11_n_351 = ~(mul_74_11_n_319 | mul_74_11_n_307);
 assign mul_74_11_n_343 = ~(mul_74_11_n_330 & ~mul_74_11_n_293);
 assign mul_74_11_n_341 = ~(mul_74_11_n_6 & n_1528);
 assign mul_74_11_n_340 = (mul_74_11_n_311 & n_1292);
 assign mul_74_11_n_339 = ~(mul_74_11_n_273 & mul_74_11_n_84);
 assign mul_74_11_n_336 = ~(mul_74_11_n_275 & mul_74_11_n_218);
 assign mul_74_11_n_335 = ~(mul_74_11_n_279 & mul_74_11_n_217);
 assign mul_74_11_n_334 = ~(mul_74_11_n_279 | mul_74_11_n_217);
 assign mul_74_11_n_333 = ~(mul_74_11_n_276 & ~mul_74_11_n_218);
 assign mul_74_11_n_332 = ~(mul_74_11_n_278 | n_1292);
 assign mul_74_11_n_331 = ~(mul_74_11_n_278 & n_1292);
 assign mul_74_11_n_330 = ~(mul_74_11_n_6 & n_1523);
 assign mul_74_11_n_342 = ~(mul_74_11_n_242 | ~mul_74_11_n_283);
 assign mul_74_11_n_328 = ~mul_74_11_n_327;
 assign mul_74_11_n_322 = ~mul_74_11_n_321;
 assign mul_74_11_n_320 = ~(mul_74_11_n_6 & n_1530);
 assign mul_74_11_n_319 = ~(mul_74_11_n_309 | mul_74_11_n_139);
 assign mul_74_11_n_318 = ~(mul_74_11_n_301 & ~(mul_74_11_n_181 & n_1487));
 assign mul_74_11_n_329 = ~(mul_74_11_n_300 | ~mul_74_11_n_205);
 assign mul_74_11_n_327 = ~(mul_74_11_n_299 | mul_74_11_n_98);
 assign mul_74_11_n_326 = ~(mul_74_11_n_302 | (mul_74_11_n_179 & n_1487));
 assign mul_74_11_n_317 = ~(mul_74_11_n_303 & (n_1514 | mul_74_11_n_47));
 assign mul_74_11_n_325 = ~(mul_74_11_n_306 | mul_74_11_n_206);
 assign mul_74_11_n_316 = ~(mul_74_11_n_304 & mul_74_11_n_207);
 assign mul_74_11_n_324 = ~(mul_74_11_n_294 & (mul_74_11_n_232 | n_1521));
 assign mul_74_11_n_323 = ~(mul_74_11_n_305 & (n_1515 | mul_74_11_n_47));
 assign mul_74_11_n_321 = ~(mul_74_11_n_297 | mul_74_11_n_208);
 assign mul_74_11_n_315 = ~(mul_74_11_n_298 & (mul_74_11_n_159 | mul_74_11_n_47));
 assign mul_74_11_n_314 = ~mul_74_11_n_313;
 assign mul_74_11_n_308 = ~(mul_74_11_n_239 & n_1528);
 assign mul_74_11_n_307 = ~(mul_74_11_n_240 | mul_74_11_n_133);
 assign mul_74_11_n_306 = ~(n_1515 | ~mul_74_11_n_255);
 assign mul_74_11_n_305 = ~(mul_74_11_n_255 & (mul_74_11_n_88 | mul_74_11_n_85));
 assign mul_74_11_n_304 = ~(mul_74_11_n_255 & (mul_74_11_n_87 | mul_74_11_n_125));
 assign mul_74_11_n_303 = ~(mul_74_11_n_255 & mul_74_11_n_181);
 assign mul_74_11_n_302 = ~(n_1514 | ~mul_74_11_n_255);
 assign mul_74_11_n_301 = ~(mul_74_11_n_255 & mul_74_11_n_180);
 assign mul_74_11_n_300 = ~(n_1506 | n_1519);
 assign mul_74_11_n_299 = ~(n_1516 | ~mul_74_11_n_255);
 assign mul_74_11_n_298 = ~(mul_74_11_n_179 & ~n_1506);
 assign mul_74_11_n_297 = ~(n_1513 | ~mul_74_11_n_255);
 assign mul_74_11_n_296 = ~(mul_74_11_n_239 & n_1530);
 assign mul_74_11_n_295 = ~(mul_74_11_n_239 & mul_74_11_n_138);
 assign mul_74_11_n_294 = ~(mul_74_11_n_239 & n_1523);
 assign mul_74_11_n_293 = ~(mul_74_11_n_240 | mul_74_11_n_139);
 assign mul_74_11_n_292 = ~(mul_74_11_n_219 | (mul_74_11_n_216 & mul_74_11_n_36));
 assign mul_74_11_n_313 = ~(mul_74_11_n_239 & n_1286);
 assign mul_74_11_n_312 = ~(mul_74_11_n_236 & mul_74_11_n_209);
 assign mul_74_11_n_291 = ~(mul_74_11_n_220 & ~(mul_74_11_n_213 & mul_74_11_n_141));
 assign mul_74_11_n_290 = ~(mul_74_11_n_221 | (n_1508 & n_1482));
 assign mul_74_11_n_289 = ~(mul_74_11_n_240 | mul_74_11_n_46);
 assign mul_74_11_n_311 = ~(mul_74_11_n_220 & ~(mul_74_11_n_213 & mul_74_11_n_31));
 assign mul_74_11_n_310 = ~(mul_74_11_n_219 | (mul_74_11_n_216 & mul_74_11_n_174));
 assign mul_74_11_n_309 = ~(mul_74_11_n_240 & mul_74_11_n_186);
 assign mul_74_11_n_287 = ~mul_74_11_n_286;
 assign mul_74_11_n_282 = ~mul_74_11_n_281;
 assign mul_74_11_n_278 = ~mul_74_11_n_277;
 assign mul_74_11_n_275 = ~mul_74_11_n_276;
 assign mul_74_11_n_273 = ~mul_74_11_n_272;
 assign mul_74_11_n_271 = ~mul_74_11_n_270;
 assign mul_74_11_n_269 = ~(mul_74_11_n_194 & ~(mul_74_11_n_213 & mul_74_11_n_128));
 assign mul_74_11_n_268 = ~((mul_74_11_n_33 | mul_74_11_n_146) & (mul_74_11_n_167 | n_1525));
 assign mul_74_11_n_267 = ~(mul_74_11_n_233 & mul_74_11_n_252);
 assign mul_74_11_n_266 = ~((mul_74_11_n_215 | mul_74_11_n_177) & (mul_74_11_n_171 | mul_74_11_n_178));
 assign mul_74_11_n_265 = ((mul_74_11_n_170 & mul_74_11_n_174) | (mul_74_11_n_216 & mul_74_11_n_223));
 assign mul_74_11_n_288 = ~(mul_74_11_n_7 | ~(mul_74_11_n_169 | n_1517));
 assign mul_74_11_n_286 = ~(mul_74_11_n_251 & ~(mul_74_11_n_216 & mul_74_11_n_176));
 assign mul_74_11_n_264 = ~((mul_74_11_n_215 | mul_74_11_n_229) & (mul_74_11_n_171 | mul_74_11_n_177));
 assign mul_74_11_n_285 = ~(mul_74_11_n_234 | mul_74_11_n_248);
 assign mul_74_11_n_284 = ~(mul_74_11_n_193 | ~mul_74_11_n_254);
 assign mul_74_11_n_283 = ~(mul_74_11_n_244 & mul_74_11_n_192);
 assign mul_74_11_n_281 = ~(mul_74_11_n_250 & ~(mul_74_11_n_216 & mul_74_11_n_225));
 assign mul_74_11_n_263 = ~(mul_74_11_n_191 & ~(n_1508 & mul_74_11_n_173));
 assign mul_74_11_n_262 = ~(mul_74_11_n_198 & ~(n_1508 & n_1520));
 assign mul_74_11_n_261 = ~(mul_74_11_n_238 & mul_74_11_n_200);
 assign mul_74_11_n_280 = ~(mul_74_11_n_235 & mul_74_11_n_199);
 assign mul_74_11_n_260 = ~(mul_74_11_n_201 & ~(n_1508 & n_1532));
 assign mul_74_11_n_279 = ~(mul_74_11_n_249 & mul_74_11_n_196);
 assign mul_74_11_n_259 = ~(mul_74_11_n_5 & ~(n_1508 & mul_74_11_n_134));
 assign mul_74_11_n_277 = ~(mul_74_11_n_246 | mul_74_11_n_195);
 assign mul_74_11_n_276 = ~(mul_74_11_n_245 | mul_74_11_n_197);
 assign mul_74_11_n_274 = ~(mul_74_11_n_237 & mul_74_11_n_202);
 assign mul_74_11_n_258 = ~(mul_74_11_n_247 & ~(n_1518 & mul_74_11_n_157));
 assign mul_74_11_n_257 = ~(mul_74_11_n_253 & ~(mul_74_11_n_216 & mul_74_11_n_222));
 assign mul_74_11_n_272 = ~(mul_74_11_n_243 | mul_74_11_n_203);
 assign mul_74_11_n_270 = ~((mul_74_11_n_216 & mul_74_11_n_224) | (mul_74_11_n_170 & mul_74_11_n_228));
 assign mul_74_11_n_255 = ~n_1506;
 assign mul_74_11_n_254 = ~(n_1510 & mul_74_11_n_157);
 assign mul_74_11_n_253 = ~(mul_74_11_n_170 & mul_74_11_n_225);
 assign mul_74_11_n_252 = ~(mul_74_11_n_170 & mul_74_11_n_222);
 assign mul_74_11_n_251 = ~(mul_74_11_n_170 & ~mul_74_11_n_175);
 assign mul_74_11_n_250 = ~(mul_74_11_n_170 & mul_74_11_n_224);
 assign mul_74_11_n_249 = ~(mul_74_11_n_213 & (mul_74_11_n_86 | mul_74_11_n_89));
 assign mul_74_11_n_248 = ~(mul_74_11_n_171 | ~mul_74_11_n_176);
 assign mul_74_11_n_247 = ~(n_1510 & n_1531);
 assign mul_74_11_n_246 = ~(n_1524 | ~mul_74_11_n_213);
 assign mul_74_11_n_245 = (mul_74_11_n_213 & n_1522);
 assign mul_74_11_n_244 = ~(n_1510 & ~n_1527);
 assign mul_74_11_n_243 = ~(n_1525 | ~n_1510);
 assign mul_74_11_n_239 = ~mul_74_11_n_240;
 assign mul_74_11_n_238 = ~(n_1508 & n_1512);
 assign mul_74_11_n_237 = ~(n_1508 & n_1534);
 assign mul_74_11_n_236 = ~(n_1508 & n_1526);
 assign mul_74_11_n_235 = ~(n_1508 & n_1533);
 assign mul_74_11_n_234 = ~(mul_74_11_n_215 | mul_74_11_n_130);
 assign mul_74_11_n_233 = ~(mul_74_11_n_216 & ~mul_74_11_n_175);
 assign mul_74_11_n_232 = ~(mul_74_11_n_166 & mul_74_11_n_186);
 assign mul_74_11_n_242 = ~(mul_74_11_n_160 & (n_1482 & mul_74_11_n_122));
 assign mul_74_11_n_231 = ~(mul_74_11_n_164 | (mul_74_11_n_30 | mul_74_11_n_119));
 assign mul_74_11_n_241 = ~(mul_74_11_n_163 | (mul_74_11_n_45 | mul_74_11_n_120));
 assign mul_74_11_n_230 = ~(mul_74_11_n_165 | (mul_74_11_n_121 | ~n_1284));
 assign mul_74_11_n_240 = ~(mul_74_11_n_102 | mul_74_11_n_101);
 assign mul_74_11_n_229 = ~mul_74_11_n_228;
 assign mul_74_11_n_227 = ~mul_74_11_n_226;
 assign mul_74_11_n_223 = ~mul_74_11_n_178;
 assign mul_74_11_n_215 = ~mul_74_11_n_216;
 assign mul_74_11_n_213 = ~mul_74_11_n_33;
 assign mul_74_11_n_33 = ~n_1510;
 assign mul_74_11_n_226 = (mul_74_11_n_36 & n_1277);
 assign mul_74_11_n_228 = (mul_74_11_n_36 ^ n_1277);
 assign mul_74_11_n_212 = (mul_74_11_n_36 & n_1279);
 assign mul_74_11_n_225 = (mul_74_11_n_36 ^ n_1279);
 assign mul_74_11_n_211 = (mul_74_11_n_36 & n_1278);
 assign mul_74_11_n_224 = (mul_74_11_n_36 ^ n_1278);
 assign mul_74_11_n_210 = (mul_74_11_n_36 & n_1280);
 assign mul_74_11_n_222 = (mul_74_11_n_36 ^ n_1280);
 assign mul_74_11_n_209 = ~(n_1512 & ~mul_74_11_n_169);
 assign mul_74_11_n_208 = ~(n_1516 | mul_74_11_n_47);
 assign mul_74_11_n_207 = ~(n_1487 & (mul_74_11_n_88 | mul_74_11_n_85));
 assign mul_74_11_n_206 = ~(n_1513 | mul_74_11_n_47);
 assign mul_74_11_n_205 = ~(mul_74_11_n_180 & n_1487);
 assign mul_74_11_n_221 = ~(mul_74_11_n_169 | mul_74_11_n_37);
 assign mul_74_11_n_220 = ~(n_1518 & mul_74_11_n_31);
 assign mul_74_11_n_204 = ~(mul_74_11_n_167 | mul_74_11_n_46);
 assign mul_74_11_n_219 = ~(mul_74_11_n_171 | mul_74_11_n_29);
 assign mul_74_11_n_218 = ~(mul_74_11_n_169 | mul_74_11_n_46);
 assign mul_74_11_n_217 = ~(mul_74_11_n_171 | mul_74_11_n_46);
 assign mul_74_11_n_216 = ~(mul_74_11_n_170 | mul_74_11_n_162);
 assign mul_74_11_n_203 = ~(n_1524 | ~n_1518);
 assign mul_74_11_n_202 = ~(n_1511 & ~mul_74_11_n_169);
 assign mul_74_11_n_201 = ~(n_1534 & ~mul_74_11_n_169);
 assign mul_74_11_n_200 = ~(n_1532 & ~mul_74_11_n_169);
 assign mul_74_11_n_199 = ~(n_1526 & ~mul_74_11_n_169);
 assign mul_74_11_n_198 = ~(n_1533 & ~mul_74_11_n_169);
 assign mul_74_11_n_197 = ~(mul_74_11_n_167 | n_1527);
 assign mul_74_11_n_196 = ~(n_1529 & ~mul_74_11_n_167);
 assign mul_74_11_n_195 = ~(mul_74_11_n_140 | ~n_1518);
 assign mul_74_11_n_194 = ~(n_1522 & ~mul_74_11_n_167);
 assign mul_74_11_n_193 = ~(mul_74_11_n_126 | ~n_1518);
 assign mul_74_11_n_192 = ~(n_1531 & ~mul_74_11_n_167);
 assign mul_74_11_n_191 = ~(mul_74_11_n_134 & ~mul_74_11_n_169);
 assign mul_74_11_n_173 = ~n_1517;
 assign mul_74_11_n_170 = ~mul_74_11_n_171;
 assign mul_74_11_n_167 = ~n_1518;
 assign mul_74_11_n_166 = ~((n_1482 & ~n_1287) | (mul_74_11_n_37 & n_1287));
 assign mul_74_11_n_165 = ~(mul_74_11_n_45 | ~(n_1285 | n_1283));
 assign mul_74_11_n_164 = ~(mul_74_11_n_117 | mul_74_11_n_35);
 assign mul_74_11_n_163 = ~(mul_74_11_n_118 | mul_74_11_n_37);
 assign mul_74_11_n_162 = ~(mul_74_11_n_110 | mul_74_11_n_0);
 assign mul_74_11_n_160 = ~(mul_74_11_n_31 & (n_1483 | n_1283));
 assign mul_74_11_n_189 = ~((n_1482 | mul_74_11_n_51) & (n_1274 | mul_74_11_n_37));
 assign mul_74_11_n_186 = ~(mul_74_11_n_99 & mul_74_11_n_100);
 assign mul_74_11_n_159 = ~(mul_74_11_n_87 | mul_74_11_n_125);
 assign mul_74_11_n_184 = ~(n_1292 & ~n_1313);
 assign mul_74_11_n_181 = ~((mul_74_11_n_35 & ~n_1479) | (n_1292 & n_1479));
 assign mul_74_11_n_180 = ~((mul_74_11_n_48 & ~n_1292) | (n_1282 & n_1292));
 assign mul_74_11_n_179 = (n_1279 ^ n_1292);
 assign mul_74_11_n_178 = ~((mul_74_11_n_29 & n_1275) | (mul_74_11_n_39 & mul_74_11_n_36));
 assign mul_74_11_n_177 = ~((mul_74_11_n_29 & n_1276) | (mul_74_11_n_50 & mul_74_11_n_36));
 assign mul_74_11_n_176 = ~((mul_74_11_n_48 & ~mul_74_11_n_36) | (n_1282 & mul_74_11_n_36));
 assign mul_74_11_n_175 = ~((n_1479 & ~mul_74_11_n_36) | (mul_74_11_n_42 & mul_74_11_n_36));
 assign mul_74_11_n_174 = ~((mul_74_11_n_36 | mul_74_11_n_51) & (n_1274 | mul_74_11_n_29));
 assign mul_74_11_n_171 = ~(mul_74_11_n_115 | mul_74_11_n_108);
 assign mul_74_11_n_169 = ~(mul_74_11_n_2 | mul_74_11_n_109);
 assign mul_74_11_n_156 = ~mul_74_11_n_155;
 assign mul_74_11_n_154 = ~mul_74_11_n_153;
 assign mul_74_11_n_146 = ~n_1529;
 assign mul_74_11_n_141 = ~mul_74_11_n_140;
 assign mul_74_11_n_130 = ~(mul_74_11_n_53 | ~(n_1283 | mul_74_11_n_29));
 assign mul_74_11_n_128 = ~((mul_74_11_n_46 & ~mul_74_11_n_31) | (n_1283 & mul_74_11_n_31));
 assign mul_74_11_n_157 = ~((mul_74_11_n_30 & ~n_1279) | (mul_74_11_n_31 & n_1279));
 assign mul_74_11_n_155 = ~((n_1286 | mul_74_11_n_41) & (n_1277 | mul_74_11_n_45));
 assign mul_74_11_n_153 = ~((mul_74_11_n_45 & n_1275) | (mul_74_11_n_39 & n_1286));
 assign mul_74_11_n_126 = ~(mul_74_11_n_86 | mul_74_11_n_89);
 assign mul_74_11_n_143 = ~((mul_74_11_n_45 & n_1276) | (mul_74_11_n_50 & n_1286));
 assign mul_74_11_n_140 = (n_1274 ^ mul_74_11_n_30);
 assign mul_74_11_n_139 = ~(mul_74_11_n_68 | ~(n_1479 | mul_74_11_n_45));
 assign mul_74_11_n_138 = ~((n_1286 | mul_74_11_n_51) & (n_1274 | mul_74_11_n_45));
 assign mul_74_11_n_134 = ~((mul_74_11_n_37 & ~n_1275) | (n_1482 & n_1275));
 assign mul_74_11_n_133 = ~(mul_74_11_n_78 | ~(n_1280 | mul_74_11_n_45));
 assign n_1313 = ~mul_74_11_n_123;
 assign mul_74_11_n_122 = ~(n_1483 & n_1283);
 assign mul_74_11_n_121 = (n_1285 & n_1283);
 assign mul_74_11_n_120 = ~(mul_74_11_n_52 | mul_74_11_n_46);
 assign mul_74_11_n_119 = (n_1486 & n_1283);
 assign mul_74_11_n_118 = ~(n_1287 | n_1283);
 assign mul_74_11_n_117 = ~(n_1486 | n_1283);
 assign mul_74_11_n_115 = ~(n_1286 | mul_74_11_n_43);
 assign mul_74_11_n_110 = ~(n_1285 | mul_74_11_n_29);
 assign mul_74_11_n_109 = ~(n_1483 | mul_74_11_n_30);
 assign mul_74_11_n_108 = ~(n_1285 | mul_74_11_n_45);
 assign mul_74_11_n_125 = ~(n_1278 | mul_74_11_n_35);
 assign mul_74_11_n_102 = ~(n_1482 | mul_74_11_n_52);
 assign mul_74_11_n_101 = ~(n_1287 | mul_74_11_n_37);
 assign mul_74_11_n_100 = ~(mul_74_11_n_45 & n_1287);
 assign mul_74_11_n_99 = ~(mul_74_11_n_52 & n_1286);
 assign mul_74_11_n_98 = ~(mul_74_11_n_47 | mul_74_11_n_35);
 assign mul_74_11_n_123 = ~(n_1487 & n_1283);
 assign mul_74_11_n_94 = ~(mul_74_11_n_36 & n_1274);
 assign mul_74_11_n_93 = ~(mul_74_11_n_29 | mul_74_11_n_39);
 assign mul_74_11_n_92 = ~(mul_74_11_n_29 | mul_74_11_n_50);
 assign mul_74_11_n_91 = ~(mul_74_11_n_29 | mul_74_11_n_42);
 assign mul_74_11_n_90 = ~(mul_74_11_n_29 | mul_74_11_n_48);
 assign mul_74_11_n_78 = ~(n_1286 | mul_74_11_n_40);
 assign mul_74_11_n_89 = ~(n_1278 | mul_74_11_n_30);
 assign mul_74_11_n_88 = ~(mul_74_11_n_41 | ~mul_74_11_n_35);
 assign mul_74_11_n_87 = ~(mul_74_11_n_38 | ~mul_74_11_n_35);
 assign mul_74_11_n_68 = ~(n_1286 | mul_74_11_n_42);
 assign mul_74_11_n_86 = ~(mul_74_11_n_38 | ~mul_74_11_n_30);
 assign mul_74_11_n_85 = ~(n_1277 | mul_74_11_n_35);
 assign mul_74_11_n_53 = ~(mul_74_11_n_36 | mul_74_11_n_46);
 assign mul_74_11_n_84 = (mul_74_11_n_36 & n_1283);
 assign mul_74_11_n_52 = ~n_1287;
 assign mul_74_11_n_51 = ~n_1274;
 assign mul_74_11_n_50 = ~n_1276;
 assign mul_74_11_n_49 = ~n_1279;
 assign mul_74_11_n_48 = ~n_1282;
 assign mul_74_11_n_47 = ~n_1487;
 assign mul_74_11_n_46 = ~n_1283;
 assign mul_74_11_n_31 = ~mul_74_11_n_30;
 assign mul_74_11_n_30 = ~n_1484;
 assign mul_74_11_n_45 = ~n_1286;
 assign mul_74_11_n_44 = ~n_1483;
 assign mul_74_11_n_43 = ~n_1285;
 assign mul_74_11_n_42 = ~n_1479;
 assign mul_74_11_n_41 = ~n_1277;
 assign mul_74_11_n_40 = ~n_1280;
 assign mul_74_11_n_39 = ~n_1275;
 assign mul_74_11_n_38 = ~n_1278;
 assign mul_74_11_n_37 = ~n_1482;
 assign mul_74_11_n_36 = ~mul_74_11_n_29;
 assign mul_74_11_n_29 = ~n_1284;
 assign mul_74_11_n_35 = ~n_1292;
 assign mul_74_11_n_27 = (mul_74_11_n_440 | mul_74_11_n_417);
 assign mul_74_11_n_26 = ~(mul_74_11_n_433 & ~mul_74_11_n_458);
 assign mul_74_11_n_25 = ~(mul_74_11_n_464 & ~mul_74_11_n_451);
 assign mul_74_11_n_24 = (mul_74_11_n_20 ^ mul_74_11_n_402);
 assign mul_74_11_n_23 = ~(mul_74_11_n_428 ^ mul_74_11_n_422);
 assign mul_74_11_n_22 = ~(mul_74_11_n_376 | ~mul_74_11_n_399);
 assign mul_74_11_n_21 = ~(mul_74_11_n_395 & ~mul_74_11_n_381);
 assign mul_74_11_n_20 = (mul_74_11_n_382 ^ mul_74_11_n_372);
 assign mul_74_11_n_19 = ~(mul_74_11_n_397 ^ n_1505);
 assign mul_74_11_n_18 = ~(mul_74_11_n_324 ^ mul_74_11_n_323);
 assign mul_74_11_n_17 = (mul_74_11_n_18 ^ mul_74_11_n_312);
 assign mul_74_11_n_16 = (mul_74_11_n_356 ^ mul_74_11_n_288);
 assign mul_74_11_n_15 = ~(mul_74_11_n_373 ^ mul_74_11_n_285);
 assign mul_74_11_n_14 = ~(mul_74_11_n_242 ^ mul_74_11_n_283);
 assign mul_74_11_n_13 = ~(mul_74_11_n_371 | ~mul_74_11_n_280);
 assign mul_74_11_n_12 = (mul_74_11_n_217 ^ mul_74_11_n_279);
 assign mul_74_11_n_11 = (mul_74_11_n_353 ^ mul_74_11_n_274);
 assign mul_74_11_n_10 = ~(mul_74_11_n_284 | ~mul_74_11_n_241);
 assign mul_74_11_n_9 = (mul_74_11_n_272 ^ mul_74_11_n_84);
 assign mul_74_11_n_8 = (mul_74_11_n_221 | (n_1508 & mul_74_11_n_189));
 assign mul_74_11_n_7 = (n_1508 & n_1511);
 assign mul_74_11_n_6 = ~(mul_74_11_n_239 | ~mul_74_11_n_186);
 assign mul_74_11_n_5 = ~(mul_74_11_n_189 & ~mul_74_11_n_169);
 assign mul_74_11_n_4 = ~(mul_74_11_n_6 & ~mul_74_11_n_133);
 assign mul_74_11_n_2 = ~(mul_74_11_n_44 | n_1484);
 assign mul_74_11_n_0 = ~(mul_74_11_n_43 | n_1284);
 assign mul_74_11_n_34 = (n_1504 ^ (mul_74_11_n_276 ^ mul_74_11_n_378));
 assign {out1[16]} = (mul_109_11_n_1217 ^ mul_109_11_n_1171);
 assign {out1[31]} = ~(mul_109_11_n_1304 ^ mul_109_11_n_1273);
 assign mul_109_11_n_1304 = ((mul_109_11_n_1303 & mul_109_11_n_1232) | ((mul_109_11_n_1232 & mul_109_11_n_1256)
    | (mul_109_11_n_1256 & mul_109_11_n_1303)));
 assign {out1[30]} = (mul_109_11_n_1232 ^ (mul_109_11_n_1256 ^ mul_109_11_n_1303));
 assign mul_109_11_n_1303 = ~(mul_109_11_n_1249 & (mul_109_11_n_1300 | mul_109_11_n_1258));
 assign {out1[29]} = ~(mul_109_11_n_1301 ^ mul_109_11_n_1267);
 assign mul_109_11_n_1301 = ~(mul_109_11_n_1248 & (mul_109_11_n_1247 | mul_109_11_n_1296));
 assign mul_109_11_n_1300 = (mul_109_11_n_1248 & (mul_109_11_n_1247 | mul_109_11_n_1296));
 assign {out1[28]} = ~(mul_109_11_n_1296 ^ mul_109_11_n_1268);
 assign {out1[27]} = ~(mul_109_11_n_1297 ^ mul_109_11_n_1269);
 assign mul_109_11_n_1297 = ~(mul_109_11_n_1265 & (mul_109_11_n_1270 | mul_109_11_n_1292));
 assign mul_109_11_n_1296 = ~(mul_109_11_n_1294 | (mul_109_11_n_1277 | (mul_109_11_n_1282 & mul_109_11_n_1278)));
 assign {out1[26]} = ~(mul_109_11_n_1292 ^ mul_109_11_n_1280);
 assign mul_109_11_n_1294 = ~(mul_109_11_n_1251 & ~(mul_109_11_n_1278 & mul_109_11_n_1290));
 assign {out1[25]} = ~(mul_109_11_n_1291 ^ mul_109_11_n_1279);
 assign mul_109_11_n_1292 = ~(mul_109_11_n_1282 | mul_109_11_n_1290);
 assign mul_109_11_n_1291 = ~(mul_109_11_n_1236 & (mul_109_11_n_1237 | mul_109_11_n_1287));
 assign mul_109_11_n_1290 = ~(mul_109_11_n_1237 | (mul_109_11_n_1287 | mul_109_11_n_1264));
 assign {out1[24]} = ~(mul_109_11_n_1287 ^ mul_109_11_n_1253);
 assign {out1[23]} = ~(mul_109_11_n_1252 ^ mul_109_11_n_1286);
 assign mul_109_11_n_1287 = ~(mul_109_11_n_1285 | ~(mul_109_11_n_1240 | mul_109_11_n_1271));
 assign mul_109_11_n_1286 = ~(mul_109_11_n_1222 & (mul_109_11_n_1276 | mul_109_11_n_1218));
 assign mul_109_11_n_1285 = ~(mul_109_11_n_1241 & (mul_109_11_n_1274 & (mul_109_11_n_1209 | mul_109_11_n_1271)));
 assign {out1[22]} = ~(mul_109_11_n_1276 ^ mul_109_11_n_1229);
 assign {out1[21]} = ~(mul_109_11_n_1275 ^ mul_109_11_n_1221);
 assign mul_109_11_n_1282 = ~(mul_109_11_n_1266 & (mul_109_11_n_1236 | mul_109_11_n_1264));
 assign {out1[19]} = ~(mul_109_11_n_1197 ^ mul_109_11_n_1261);
 assign mul_109_11_n_1280 = ~(mul_109_11_n_1270 | ~mul_109_11_n_1265);
 assign mul_109_11_n_1279 = ~(mul_109_11_n_1266 & ~mul_109_11_n_1264);
 assign mul_109_11_n_1278 = ~(mul_109_11_n_1270 | mul_109_11_n_1246);
 assign mul_109_11_n_1277 = ~(mul_109_11_n_1265 | mul_109_11_n_1246);
 assign mul_109_11_n_1276 = ~(mul_109_11_n_1228 | (mul_109_11_n_1219 & mul_109_11_n_1257));
 assign mul_109_11_n_1275 = ~(mul_109_11_n_1212 & ~(mul_109_11_n_1210 & mul_109_11_n_1257));
 assign mul_109_11_n_1274 = ~(mul_109_11_n_1254 | (mul_109_11_n_1228 & mul_109_11_n_1250));
 assign mul_109_11_n_1273 = ~(mul_109_11_n_1234 ^ mul_109_11_n_1255);
 assign {out1[20]} = ~(mul_109_11_n_1257 ^ mul_109_11_n_1220);
 assign mul_109_11_n_1269 = ~(mul_109_11_n_1251 & ~mul_109_11_n_1246);
 assign mul_109_11_n_1268 = ~(mul_109_11_n_1247 | ~mul_109_11_n_1248);
 assign mul_109_11_n_1267 = ~(mul_109_11_n_1249 & ~mul_109_11_n_1258);
 assign mul_109_11_n_1271 = ~(mul_109_11_n_1250 & mul_109_11_n_1219);
 assign mul_109_11_n_1270 = ~(mul_109_11_n_1259 | mul_109_11_n_1226);
 assign {out1[18]} = ~(mul_109_11_n_1187 ^ mul_109_11_n_1239);
 assign {out1[17]} = ~(mul_109_11_n_1235 ^ mul_109_11_n_1170);
 assign mul_109_11_n_1266 = ~(mul_109_11_n_1260 & mul_109_11_n_1223);
 assign mul_109_11_n_1261 = ~(mul_109_11_n_1177 & (mul_109_11_n_1168 | mul_109_11_n_1239));
 assign mul_109_11_n_1265 = ~(mul_109_11_n_1259 & mul_109_11_n_1226);
 assign mul_109_11_n_1264 = ~(mul_109_11_n_1260 | mul_109_11_n_1223);
 assign mul_109_11_n_1259 = ((mul_109_11_n_1146 & mul_109_11_n_1202) | ((mul_109_11_n_1202 & mul_109_11_n_1131)
    | (mul_109_11_n_1131 & mul_109_11_n_1146)));
 assign mul_109_11_n_1260 = (mul_109_11_n_1202 ^ (mul_109_11_n_1131 ^ mul_109_11_n_1146));
 assign mul_109_11_n_1255 = ((mul_109_11_n_1208 & mul_109_11_n_1140) | ((mul_109_11_n_1140 & mul_109_11_n_1198)
    | (mul_109_11_n_1198 & mul_109_11_n_1208)));
 assign mul_109_11_n_1256 = (mul_109_11_n_1140 ^ (mul_109_11_n_1198 ^ mul_109_11_n_1208));
 assign mul_109_11_n_1254 = ~(mul_109_11_n_1238 | mul_109_11_n_1222);
 assign mul_109_11_n_1253 = ~(mul_109_11_n_1237 | ~mul_109_11_n_1236);
 assign mul_109_11_n_1252 = ~(mul_109_11_n_1241 & ~mul_109_11_n_1238);
 assign mul_109_11_n_1258 = ~(mul_109_11_n_1244 | mul_109_11_n_1233);
 assign mul_109_11_n_1257 = ~(mul_109_11_n_1209 & mul_109_11_n_1240);
 assign mul_109_11_n_1251 = ~(mul_109_11_n_1243 & mul_109_11_n_1225);
 assign mul_109_11_n_1250 = ~(mul_109_11_n_1238 | mul_109_11_n_1218);
 assign mul_109_11_n_1249 = ~(mul_109_11_n_1244 & mul_109_11_n_1233);
 assign mul_109_11_n_1248 = ~(mul_109_11_n_1242 & mul_109_11_n_1245);
 assign mul_109_11_n_1247 = ~(mul_109_11_n_1242 | mul_109_11_n_1245);
 assign mul_109_11_n_1246 = ~(mul_109_11_n_1243 | mul_109_11_n_1225);
 assign mul_109_11_n_1244 = ((mul_109_11_n_1176 & mul_109_11_n_1190) | ((mul_109_11_n_1190 & mul_109_11_n_1133)
    | (mul_109_11_n_1133 & mul_109_11_n_1176)));
 assign mul_109_11_n_1245 = (mul_109_11_n_1190 ^ (mul_109_11_n_1133 ^ mul_109_11_n_1176));
 assign mul_109_11_n_1242 = ((mul_109_11_n_1191 & mul_109_11_n_1188) | ((mul_109_11_n_1188 & mul_109_11_n_1115)
    | (mul_109_11_n_1115 & mul_109_11_n_1191)));
 assign mul_109_11_n_1243 = (mul_109_11_n_1188 ^ (mul_109_11_n_1115 ^ mul_109_11_n_1191));
 assign mul_109_11_n_1241 = ~(mul_109_11_n_1231 & mul_109_11_n_1214);
 assign mul_109_11_n_1240 = ~(mul_109_11_n_1227 & mul_109_11_n_1195);
 assign mul_109_11_n_1239 = ~(mul_109_11_n_1227 | mul_109_11_n_1182);
 assign mul_109_11_n_1238 = ~(mul_109_11_n_1231 | mul_109_11_n_1214);
 assign mul_109_11_n_1235 = ~(mul_109_11_n_1158 & (mul_109_11_n_1160 | mul_109_11_n_1217));
 assign mul_109_11_n_1234 = ~(mul_109_11_n_1165 ^ mul_109_11_n_1216);
 assign mul_109_11_n_1237 = ~(mul_109_11_n_1230 | mul_109_11_n_1224);
 assign mul_109_11_n_1236 = ~(mul_109_11_n_1230 & mul_109_11_n_1224);
 assign mul_109_11_n_1232 = ((mul_109_11_n_1199 & mul_109_11_n_1175) | ((mul_109_11_n_1175 & mul_109_11_n_1157)
    | (mul_109_11_n_1157 & mul_109_11_n_1199)));
 assign mul_109_11_n_1233 = (mul_109_11_n_1175 ^ (mul_109_11_n_1157 ^ mul_109_11_n_1199));
 assign mul_109_11_n_1230 = ((mul_109_11_n_1129 & mul_109_11_n_1173) | ((mul_109_11_n_1173 & mul_109_11_n_1113)
    | (mul_109_11_n_1113 & mul_109_11_n_1129)));
 assign mul_109_11_n_1231 = (mul_109_11_n_1173 ^ (mul_109_11_n_1113 ^ mul_109_11_n_1129));
 assign mul_109_11_n_1229 = ~(mul_109_11_n_1218 | ~mul_109_11_n_1222);
 assign mul_109_11_n_1228 = ~(mul_109_11_n_1211 & (mul_109_11_n_1212 | mul_109_11_n_1213));
 assign mul_109_11_n_1227 = ~(mul_109_11_n_1160 | (mul_109_11_n_1159 | mul_109_11_n_1217));
 assign mul_109_11_n_1225 = ((mul_109_11_n_1145 & mul_109_11_n_1189) | ((mul_109_11_n_1189 & mul_109_11_n_1117)
    | (mul_109_11_n_1117 & mul_109_11_n_1145)));
 assign mul_109_11_n_1226 = (mul_109_11_n_1189 ^ (mul_109_11_n_1117 ^ mul_109_11_n_1145));
 assign mul_109_11_n_1223 = ((mul_109_11_n_1203 & mul_109_11_n_1128) | ((mul_109_11_n_1128 & mul_109_11_n_1084)
    | (mul_109_11_n_1084 & mul_109_11_n_1203)));
 assign mul_109_11_n_1224 = (mul_109_11_n_1128 ^ (mul_109_11_n_1084 ^ mul_109_11_n_1203));
 assign mul_109_11_n_1221 = ~(mul_109_11_n_1211 & ~mul_109_11_n_1213);
 assign mul_109_11_n_1220 = ~(mul_109_11_n_1210 & mul_109_11_n_1212);
 assign mul_109_11_n_1222 = ~(mul_109_11_n_1200 & mul_109_11_n_1215);
 assign mul_109_11_n_1219 = ~(mul_109_11_n_1213 | ~mul_109_11_n_1210);
 assign mul_109_11_n_1216 = ~(mul_109_11_n_1207 ^ mul_109_11_n_1166);
 assign mul_109_11_n_1218 = ~(mul_109_11_n_1200 | mul_109_11_n_1215);
 assign mul_109_11_n_1217 = ~(mul_109_11_n_1194 | (mul_109_11_n_1167 | (mul_109_11_n_1192 | mul_109_11_n_1193)));
 assign mul_109_11_n_1214 = ((mul_109_11_n_1143 & mul_109_11_n_1174) | ((mul_109_11_n_1174 & mul_109_11_n_1019)
    | (mul_109_11_n_1019 & mul_109_11_n_1143)));
 assign mul_109_11_n_1215 = (mul_109_11_n_1174 ^ (mul_109_11_n_1019 ^ mul_109_11_n_1143));
 assign mul_109_11_n_1213 = ~(mul_109_11_n_1205 | mul_109_11_n_1201);
 assign mul_109_11_n_1212 = ~(mul_109_11_n_1206 & mul_109_11_n_1178);
 assign mul_109_11_n_1211 = ~(mul_109_11_n_1205 & mul_109_11_n_1201);
 assign mul_109_11_n_1210 = (mul_109_11_n_1206 | mul_109_11_n_1178);
 assign mul_109_11_n_1209 = ~(mul_109_11_n_1196 | (mul_109_11_n_1186 | (mul_109_11_n_1195 & mul_109_11_n_1182)));
 assign mul_109_11_n_1207 = ((mul_109_11_n_1080 & mul_109_11_n_1156) | ((mul_109_11_n_1156 & mul_109_11_n_1142)
    | (mul_109_11_n_1142 & mul_109_11_n_1080)));
 assign mul_109_11_n_1208 = (mul_109_11_n_1156 ^ (mul_109_11_n_1142 ^ mul_109_11_n_1080));
 assign mul_109_11_n_1205 = ((mul_109_11_n_1111 & mul_109_11_n_1126) | ((mul_109_11_n_1126 & mul_109_11_n_1043)
    | (mul_109_11_n_1043 & mul_109_11_n_1111)));
 assign mul_109_11_n_1206 = (mul_109_11_n_1126 ^ (mul_109_11_n_1043 ^ mul_109_11_n_1111));
 assign {out1[15]} = ~(mul_109_11_n_1172 ^ mul_109_11_n_1183);
 assign mul_109_11_n_1202 = ((mul_109_11_n_1027 & mul_109_11_n_1022) | ((mul_109_11_n_1022 & mul_109_11_n_1112)
    | (mul_109_11_n_1112 & mul_109_11_n_1027)));
 assign mul_109_11_n_1203 = (mul_109_11_n_1022 ^ (mul_109_11_n_1112 ^ mul_109_11_n_1027));
 assign mul_109_11_n_1200 = ((mul_109_11_n_1144 & mul_109_11_n_1110) | ((mul_109_11_n_1110 & mul_109_11_n_1042)
    | (mul_109_11_n_1042 & mul_109_11_n_1144)));
 assign mul_109_11_n_1201 = (mul_109_11_n_1110 ^ (mul_109_11_n_1042 ^ mul_109_11_n_1144));
 assign mul_109_11_n_1198 = ((mul_109_11_n_1132 & mul_109_11_n_1100) | ((mul_109_11_n_1100 & mul_109_11_n_1081)
    | (mul_109_11_n_1081 & mul_109_11_n_1132)));
 assign mul_109_11_n_1199 = (mul_109_11_n_1100 ^ (mul_109_11_n_1081 ^ mul_109_11_n_1132));
 assign mul_109_11_n_1197 = (mul_109_11_n_1185 | mul_109_11_n_1186);
 assign mul_109_11_n_1196 = ~(mul_109_11_n_1185 | mul_109_11_n_1177);
 assign mul_109_11_n_1195 = ~(mul_109_11_n_1185 | mul_109_11_n_1168);
 assign mul_109_11_n_1194 = ~(mul_109_11_n_1184 | ~mul_109_11_n_1108);
 assign mul_109_11_n_1193 = ~(mul_109_11_n_1184 | mul_109_11_n_1093);
 assign mul_109_11_n_1192 = ~(mul_109_11_n_1155 & ~(mul_109_11_n_1169 & mul_109_11_n_1123));
 assign mul_109_11_n_1190 = ((mul_109_11_n_1116 & mul_109_11_n_1095) | ((mul_109_11_n_1095 & mul_109_11_n_1068)
    | (mul_109_11_n_1068 & mul_109_11_n_1116)));
 assign mul_109_11_n_1191 = (mul_109_11_n_1095 ^ (mul_109_11_n_1068 ^ mul_109_11_n_1116));
 assign mul_109_11_n_1188 = ((mul_109_11_n_1130 & mul_109_11_n_1009) | ((mul_109_11_n_1009 & mul_109_11_n_1096)
    | (mul_109_11_n_1096 & mul_109_11_n_1130)));
 assign mul_109_11_n_1189 = (mul_109_11_n_1009 ^ (mul_109_11_n_1096 ^ mul_109_11_n_1130));
 assign mul_109_11_n_1187 = ~(mul_109_11_n_1168 | ~mul_109_11_n_1177);
 assign mul_109_11_n_1186 = (mul_109_11_n_1163 & mul_109_11_n_1179);
 assign mul_109_11_n_1185 = ~(mul_109_11_n_1163 | mul_109_11_n_1179);
 assign mul_109_11_n_1184 = ~(mul_109_11_n_1120 & mul_109_11_n_1169);
 assign mul_109_11_n_1183 = ~(mul_109_11_n_1119 & (mul_109_11_n_1118 | mul_109_11_n_1154));
 assign mul_109_11_n_1182 = ~(mul_109_11_n_1162 & (mul_109_11_n_1158 | mul_109_11_n_1159));
 assign {out1[14]} = ~(mul_109_11_n_1125 ^ mul_109_11_n_1154);
 assign {out1[13]} = ~(mul_109_11_n_1109 ^ mul_109_11_n_1151);
 assign mul_109_11_n_1175 = ((mul_109_11_n_1114 & mul_109_11_n_1082) | ((mul_109_11_n_1082 & mul_109_11_n_1047)
    | (mul_109_11_n_1047 & mul_109_11_n_1114)));
 assign mul_109_11_n_1176 = (mul_109_11_n_1082 ^ (mul_109_11_n_1047 ^ mul_109_11_n_1114));
 assign mul_109_11_n_1178 = ((mul_109_11_n_1127 & mul_109_11_n_1041) | ((mul_109_11_n_1041 & mul_109_11_n_1085)
    | (mul_109_11_n_1085 & mul_109_11_n_1127)));
 assign mul_109_11_n_1179 = (mul_109_11_n_1041 ^ (mul_109_11_n_1085 ^ mul_109_11_n_1127));
 assign mul_109_11_n_1173 = ((mul_109_11_n_1097 & mul_109_11_n_1070) | ((mul_109_11_n_1070 & mul_109_11_n_1050)
    | (mul_109_11_n_1050 & mul_109_11_n_1097)));
 assign mul_109_11_n_1174 = (mul_109_11_n_1070 ^ (mul_109_11_n_1050 ^ mul_109_11_n_1097));
 assign mul_109_11_n_1172 = ~(mul_109_11_n_1155 & ~mul_109_11_n_1161);
 assign mul_109_11_n_1171 = ~(mul_109_11_n_1158 & ~mul_109_11_n_1160);
 assign mul_109_11_n_1170 = ~(mul_109_11_n_1162 & ~mul_109_11_n_1159);
 assign mul_109_11_n_1177 = ~(mul_109_11_n_1164 & mul_109_11_n_1149);
 assign mul_109_11_n_1167 = ~(mul_109_11_n_1161 | mul_109_11_n_1119);
 assign mul_109_11_n_1169 = ~(mul_109_11_n_1161 | mul_109_11_n_1118);
 assign mul_109_11_n_1166 = ~(mul_109_11_n_1107 ^ mul_109_11_n_1141);
 assign mul_109_11_n_1165 = ~(mul_109_11_n_1138 ^ mul_109_11_n_1139);
 assign mul_109_11_n_1168 = ~(mul_109_11_n_1164 | mul_109_11_n_1149);
 assign mul_109_11_n_1163 = ((mul_109_11_n_1086 & mul_109_11_n_1037) | ((mul_109_11_n_1037 & mul_109_11_n_1073)
    | (mul_109_11_n_1073 & mul_109_11_n_1086)));
 assign mul_109_11_n_1164 = (mul_109_11_n_1037 ^ (mul_109_11_n_1073 ^ mul_109_11_n_1086));
 assign mul_109_11_n_1156 = ((mul_109_11_n_1053 & mul_109_11_n_1046) | ((mul_109_11_n_1046 & mul_109_11_n_1072)
    | (mul_109_11_n_1072 & mul_109_11_n_1053)));
 assign mul_109_11_n_1157 = (mul_109_11_n_1046 ^ (mul_109_11_n_1072 ^ mul_109_11_n_1053));
 assign mul_109_11_n_1162 = ~(mul_109_11_n_1150 & mul_109_11_n_1136);
 assign mul_109_11_n_1161 = ~(mul_109_11_n_1148 | mul_109_11_n_1103);
 assign mul_109_11_n_1160 = ~(mul_109_11_n_1137 | mul_109_11_n_1147);
 assign mul_109_11_n_1159 = ~(mul_109_11_n_1150 | mul_109_11_n_1136);
 assign mul_109_11_n_1158 = ~(mul_109_11_n_1137 & mul_109_11_n_1147);
 assign {out1[11]} = ~(mul_109_11_n_1015 ^ mul_109_11_n_1124);
 assign {out1[12]} = ~(mul_109_11_n_1135 ^ mul_109_11_n_1078);
 assign mul_109_11_n_1155 = ~(mul_109_11_n_1148 & mul_109_11_n_1103);
 assign mul_109_11_n_1151 = ~(mul_109_11_n_1063 & (mul_109_11_n_1135 | mul_109_11_n_1064));
 assign mul_109_11_n_1154 = ~(mul_109_11_n_1123 | (mul_109_11_n_1120 & mul_109_11_n_1134));
 assign mul_109_11_n_1149 = ((mul_109_11_n_1074 & mul_109_11_n_1003) | ((mul_109_11_n_1003 & mul_109_11_n_1056)
    | (mul_109_11_n_1056 & mul_109_11_n_1074)));
 assign mul_109_11_n_1150 = (mul_109_11_n_1003 ^ (mul_109_11_n_1056 ^ mul_109_11_n_1074));
 assign mul_109_11_n_1147 = ((mul_109_11_n_1025 & mul_109_11_n_952) | ((mul_109_11_n_952 & mul_109_11_n_1054)
    | (mul_109_11_n_1054 & mul_109_11_n_1025)));
 assign mul_109_11_n_1148 = (mul_109_11_n_952 ^ (mul_109_11_n_1054 ^ mul_109_11_n_1025));
 assign mul_109_11_n_1145 = ((mul_109_11_n_1083 & mul_109_11_n_1039) | ((mul_109_11_n_1039 & mul_109_11_n_1026)
    | (mul_109_11_n_1026 & mul_109_11_n_1083)));
 assign mul_109_11_n_1146 = (mul_109_11_n_1039 ^ (mul_109_11_n_1026 ^ mul_109_11_n_1083));
 assign mul_109_11_n_1143 = ((mul_109_11_n_1098 & mul_109_11_n_737) | ((mul_109_11_n_737 & mul_109_11_n_1051)
    | (mul_109_11_n_1051 & mul_109_11_n_1098)));
 assign mul_109_11_n_1144 = (mul_109_11_n_737 ^ (mul_109_11_n_1051 ^ mul_109_11_n_1098));
 assign mul_109_11_n_1141 = ((mul_109_11_n_1071 & mul_109_11_n_639) | ((mul_109_11_n_639 & mul_109_11_n_1049)
    | (mul_109_11_n_1049 & mul_109_11_n_1071)));
 assign mul_109_11_n_1142 = (mul_109_11_n_639 ^ (mul_109_11_n_1049 ^ mul_109_11_n_1071));
 assign mul_109_11_n_1139 = ((mul_109_11_n_1099 & mul_109_11_n_1052) | ((mul_109_11_n_1052 & mul_109_11_n_1045)
    | (mul_109_11_n_1045 & mul_109_11_n_1099)));
 assign mul_109_11_n_1140 = (mul_109_11_n_1052 ^ (mul_109_11_n_1045 ^ mul_109_11_n_1099));
 assign mul_109_11_n_1138 = ~(mul_109_11_n_1105 ^ mul_109_11_n_1106);
 assign mul_109_11_n_1135 = ~mul_109_11_n_1134;
 assign mul_109_11_n_1132 = ((mul_109_11_n_1067 & mul_109_11_n_980) | ((mul_109_11_n_980 & mul_109_11_n_1028)
    | (mul_109_11_n_1028 & mul_109_11_n_1067)));
 assign mul_109_11_n_1133 = (mul_109_11_n_980 ^ (mul_109_11_n_1028 ^ mul_109_11_n_1067));
 assign mul_109_11_n_1136 = ((mul_109_11_n_1057 & mul_109_11_n_935) | ((mul_109_11_n_935 & mul_109_11_n_1024)
    | (mul_109_11_n_1024 & mul_109_11_n_1057)));
 assign mul_109_11_n_1137 = (mul_109_11_n_935 ^ (mul_109_11_n_1024 ^ mul_109_11_n_1057));
 assign mul_109_11_n_1130 = ((mul_109_11_n_960 & mul_109_11_n_1021) | ((mul_109_11_n_1021 & mul_109_11_n_1010)
    | (mul_109_11_n_1010 & mul_109_11_n_960)));
 assign mul_109_11_n_1131 = (mul_109_11_n_1021 ^ (mul_109_11_n_1010 ^ mul_109_11_n_960));
 assign mul_109_11_n_1128 = ((mul_109_11_n_1023 & mul_109_11_n_969) | ((mul_109_11_n_969 & mul_109_11_n_1018)
    | (mul_109_11_n_1018 & mul_109_11_n_1023)));
 assign mul_109_11_n_1129 = (mul_109_11_n_969 ^ (mul_109_11_n_1018 ^ mul_109_11_n_1023));
 assign mul_109_11_n_1126 = ((mul_109_11_n_1036 & mul_109_11_n_984) | ((mul_109_11_n_984 & mul_109_11_n_923)
    | (mul_109_11_n_923 & mul_109_11_n_1036)));
 assign mul_109_11_n_1127 = (mul_109_11_n_984 ^ (mul_109_11_n_923 ^ mul_109_11_n_1036));
 assign mul_109_11_n_1125 = ~(mul_109_11_n_1118 | ~mul_109_11_n_1119);
 assign mul_109_11_n_1124 = ~(mul_109_11_n_1012 & (mul_109_11_n_1102 | mul_109_11_n_998));
 assign mul_109_11_n_1134 = ~(mul_109_11_n_1093 & ~mul_109_11_n_1108);
 assign {out1[10]} = ~(mul_109_11_n_1017 ^ mul_109_11_n_1102);
 assign {out1[9]} = ~(mul_109_11_n_1066 ^ mul_109_11_n_1090);
 assign mul_109_11_n_1123 = ~(mul_109_11_n_1092 & (mul_109_11_n_1101 | mul_109_11_n_1063));
 assign mul_109_11_n_1116 = ((mul_109_11_n_967 & mul_109_11_n_1038) | ((mul_109_11_n_1038 & mul_109_11_n_959)
    | (mul_109_11_n_959 & mul_109_11_n_967)));
 assign mul_109_11_n_1117 = (mul_109_11_n_1038 ^ (mul_109_11_n_959 ^ mul_109_11_n_967));
 assign mul_109_11_n_1114 = ((mul_109_11_n_1029 & mul_109_11_n_834) | ((mul_109_11_n_834 & mul_109_11_n_1008)
    | (mul_109_11_n_1008 & mul_109_11_n_1029)));
 assign mul_109_11_n_1115 = (mul_109_11_n_834 ^ (mul_109_11_n_1008 ^ mul_109_11_n_1029));
 assign mul_109_11_n_1112 = ((mul_109_11_n_1069 & mul_109_11_n_954) | ((mul_109_11_n_954 & mul_109_11_n_906)
    | (mul_109_11_n_906 & mul_109_11_n_1069)));
 assign mul_109_11_n_1113 = (mul_109_11_n_954 ^ (mul_109_11_n_906 ^ mul_109_11_n_1069));
 assign mul_109_11_n_1110 = ((mul_109_11_n_1007 & mul_109_11_n_1040) | ((mul_109_11_n_1040 & mul_109_11_n_983)
    | (mul_109_11_n_983 & mul_109_11_n_1007)));
 assign mul_109_11_n_1111 = (mul_109_11_n_1040 ^ (mul_109_11_n_983 ^ mul_109_11_n_1007));
 assign mul_109_11_n_1120 = ~(mul_109_11_n_1101 | mul_109_11_n_1064);
 assign mul_109_11_n_1109 = ~(mul_109_11_n_1092 & ~mul_109_11_n_1101);
 assign mul_109_11_n_1119 = ~(mul_109_11_n_1104 & mul_109_11_n_1088);
 assign mul_109_11_n_1118 = ~(mul_109_11_n_1104 | mul_109_11_n_1088);
 assign mul_109_11_n_1107 = ~(mul_109_11_n_1079 ^ mul_109_11_n_1014);
 assign mul_109_11_n_1106 = ~(mul_109_11_n_1076 ^ mul_109_11_n_918);
 assign mul_109_11_n_1105 = ~(mul_109_11_n_1075 ^ mul_109_11_n_997);
 assign mul_109_11_n_1108 = ~(mul_109_11_n_1013 & (mul_109_11_n_1094 & (mul_109_11_n_999 | mul_109_11_n_1012)));
 assign mul_109_11_n_1103 = ((mul_109_11_n_1055 & mul_109_11_n_917) | ((mul_109_11_n_917 & mul_109_11_n_961)
    | (mul_109_11_n_961 & mul_109_11_n_1055)));
 assign mul_109_11_n_1104 = (mul_109_11_n_917 ^ (mul_109_11_n_961 ^ mul_109_11_n_1055));
 assign mul_109_11_n_1099 = ((mul_109_11_n_979 & mul_109_11_n_948) | ((mul_109_11_n_948 & mul_109_11_n_975)
    | (mul_109_11_n_975 & mul_109_11_n_979)));
 assign mul_109_11_n_1100 = (mul_109_11_n_948 ^ (mul_109_11_n_975 ^ mul_109_11_n_979));
 assign mul_109_11_n_1097 = ((mul_109_11_n_1005 & mul_109_11_n_505) | ((mul_109_11_n_505 & mul_109_11_n_1006)
    | (mul_109_11_n_1006 & mul_109_11_n_1005)));
 assign mul_109_11_n_1098 = (mul_109_11_n_505 ^ (mul_109_11_n_1006 ^ mul_109_11_n_1005));
 assign mul_109_11_n_1095 = ((mul_109_11_n_946 & mul_109_11_n_509) | ((mul_109_11_n_509 & mul_109_11_n_1020)
    | (mul_109_11_n_1020 & mul_109_11_n_946)));
 assign mul_109_11_n_1096 = (mul_109_11_n_509 ^ (mul_109_11_n_1020 ^ mul_109_11_n_946));
 assign mul_109_11_n_1094 = ~(mul_109_11_n_1030 & mul_109_11_n_1087);
 assign mul_109_11_n_1102 = ~(mul_109_11_n_1077 | mul_109_11_n_1087);
 assign mul_109_11_n_1101 = ~(mul_109_11_n_1089 | mul_109_11_n_1060);
 assign {out1[8]} = ~(mul_109_11_n_1065 ^ mul_109_11_n_1062);
 assign mul_109_11_n_1093 = ~(mul_109_11_n_1077 & mul_109_11_n_1030);
 assign mul_109_11_n_1092 = ~(mul_109_11_n_1089 & mul_109_11_n_1060);
 assign mul_109_11_n_1090 = ~(mul_109_11_n_1058 & (mul_109_11_n_1062 | mul_109_11_n_1035));
 assign mul_109_11_n_1085 = ((mul_109_11_n_982 & mul_109_11_n_1002) | ((mul_109_11_n_1002 & mul_109_11_n_911)
    | (mul_109_11_n_911 & mul_109_11_n_982)));
 assign mul_109_11_n_1086 = (mul_109_11_n_1002 ^ (mul_109_11_n_911 ^ mul_109_11_n_982));
 assign mul_109_11_n_1083 = ((mul_109_11_n_1011 & mul_109_11_n_958) | ((mul_109_11_n_958 & mul_109_11_n_968)
    | (mul_109_11_n_968 & mul_109_11_n_1011)));
 assign mul_109_11_n_1084 = (mul_109_11_n_958 ^ (mul_109_11_n_968 ^ mul_109_11_n_1011));
 assign mul_109_11_n_1081 = ((mul_109_11_n_976 & mul_109_11_n_833) | ((mul_109_11_n_833 & mul_109_11_n_963)
    | (mul_109_11_n_963 & mul_109_11_n_976)));
 assign mul_109_11_n_1082 = (mul_109_11_n_833 ^ (mul_109_11_n_963 ^ mul_109_11_n_976));
 assign mul_109_11_n_1088 = ((mul_109_11_n_990 & mul_109_11_n_962) | ((mul_109_11_n_962 & mul_109_11_n_949)
    | (mul_109_11_n_949 & mul_109_11_n_990)));
 assign mul_109_11_n_1089 = (mul_109_11_n_962 ^ (mul_109_11_n_949 ^ mul_109_11_n_990));
 assign mul_109_11_n_1079 = ((mul_109_11_n_986 & mul_109_11_n_947) | ((mul_109_11_n_947 & mul_109_11_n_619)
    | (mul_109_11_n_619 & mul_109_11_n_986)));
 assign mul_109_11_n_1080 = (mul_109_11_n_947 ^ (mul_109_11_n_619 ^ mul_109_11_n_986));
 assign mul_109_11_n_1078 = ~(mul_109_11_n_1064 | ~mul_109_11_n_1063);
 assign mul_109_11_n_1087 = ~(mul_109_11_n_1059 & (mul_109_11_n_1034 | mul_109_11_n_1058));
 assign mul_109_11_n_1077 = ~(mul_109_11_n_1034 | (mul_109_11_n_1035 | mul_109_11_n_1062));
 assign mul_109_11_n_1076 = ~(mul_109_11_n_679 ^ mul_109_11_n_1048);
 assign mul_109_11_n_1075 = ~(mul_109_11_n_545 ^ mul_109_11_n_1044);
 assign mul_109_11_n_1073 = ((mul_109_11_n_934 & mul_109_11_n_978) | ((mul_109_11_n_978 & mul_109_11_n_855)
    | (mul_109_11_n_855 & mul_109_11_n_934)));
 assign mul_109_11_n_1074 = (mul_109_11_n_978 ^ (mul_109_11_n_855 ^ mul_109_11_n_934));
 assign mul_109_11_n_1071 = ((mul_109_11_n_944 & mul_109_11_n_510) | ((mul_109_11_n_510 & mul_109_11_n_939)
    | (mul_109_11_n_939 & mul_109_11_n_944)));
 assign mul_109_11_n_1072 = (mul_109_11_n_510 ^ (mul_109_11_n_939 ^ mul_109_11_n_944));
 assign mul_109_11_n_1069 = ((mul_109_11_n_1004 & mul_109_11_n_504) | ((mul_109_11_n_504 & mul_109_11_n_876)
    | (mul_109_11_n_876 & mul_109_11_n_1004)));
 assign mul_109_11_n_1070 = (mul_109_11_n_504 ^ (mul_109_11_n_876 ^ mul_109_11_n_1004));
 assign mul_109_11_n_1067 = ((mul_109_11_n_966 & mul_109_11_n_668) | ((mul_109_11_n_668 & mul_109_11_n_964)
    | (mul_109_11_n_964 & mul_109_11_n_966)));
 assign mul_109_11_n_1068 = (mul_109_11_n_668 ^ (mul_109_11_n_964 ^ mul_109_11_n_966));
 assign mul_109_11_n_1066 = ~(mul_109_11_n_1059 & ~mul_109_11_n_1034);
 assign mul_109_11_n_1065 = ~(mul_109_11_n_1035 | ~mul_109_11_n_1058);
 assign mul_109_11_n_1064 = ~(mul_109_11_n_1061 | mul_109_11_n_993);
 assign mul_109_11_n_1063 = ~(mul_109_11_n_1061 & mul_109_11_n_993);
 assign mul_109_11_n_1062 = ~(mul_109_11_n_1016 | ((mul_109_11_n_1000 & mul_109_11_n_902) | (mul_109_11_n_1000
    & mul_109_11_n_936)));
 assign mul_109_11_n_1056 = ((mul_109_11_n_951 & mul_109_11_n_905) | ((mul_109_11_n_905 & mul_109_11_n_932)
    | (mul_109_11_n_932 & mul_109_11_n_951)));
 assign mul_109_11_n_1057 = (mul_109_11_n_905 ^ (mul_109_11_n_932 ^ mul_109_11_n_951));
 assign mul_109_11_n_1054 = ((mul_109_11_n_989 & mul_109_11_n_846) | ((mul_109_11_n_846 & mul_109_11_n_871)
    | (mul_109_11_n_871 & mul_109_11_n_989)));
 assign mul_109_11_n_1055 = (mul_109_11_n_846 ^ (mul_109_11_n_871 ^ mul_109_11_n_989));
 assign mul_109_11_n_1060 = ((mul_109_11_n_950 & mul_109_11_n_870) | ((mul_109_11_n_870 & mul_109_11_n_928)
    | (mul_109_11_n_928 & mul_109_11_n_950)));
 assign mul_109_11_n_1061 = (mul_109_11_n_870 ^ (mul_109_11_n_928 ^ mul_109_11_n_950));
 assign mul_109_11_n_1052 = ((mul_109_11_n_942 & mul_109_11_n_622) | ((mul_109_11_n_622 & mul_109_11_n_669)
    | (mul_109_11_n_669 & mul_109_11_n_942)));
 assign mul_109_11_n_1053 = (mul_109_11_n_622 ^ (mul_109_11_n_669 ^ mul_109_11_n_942));
 assign mul_109_11_n_1050 = ((mul_109_11_n_987 & mul_109_11_n_812) | ((mul_109_11_n_812 & mul_109_11_n_837)
    | (mul_109_11_n_837 & mul_109_11_n_987)));
 assign mul_109_11_n_1051 = (mul_109_11_n_812 ^ (mul_109_11_n_837 ^ mul_109_11_n_987));
 assign mul_109_11_n_1048 = ((mul_109_11_n_943 & mul_109_11_n_511) | ((mul_109_11_n_511 & mul_109_11_n_861)
    | (mul_109_11_n_861 & mul_109_11_n_943)));
 assign mul_109_11_n_1049 = (mul_109_11_n_511 ^ (mul_109_11_n_861 ^ mul_109_11_n_943));
 assign mul_109_11_n_1046 = ((mul_109_11_n_940 & mul_109_11_n_670) | ((mul_109_11_n_670 & mul_109_11_n_930)
    | (mul_109_11_n_930 & mul_109_11_n_940)));
 assign mul_109_11_n_1047 = (mul_109_11_n_670 ^ (mul_109_11_n_930 ^ mul_109_11_n_940));
 assign mul_109_11_n_1044 = ((mul_109_11_n_941 & mul_109_11_n_382) | ((mul_109_11_n_382 & mul_109_11_n_925)
    | (mul_109_11_n_925 & mul_109_11_n_941)));
 assign mul_109_11_n_1045 = (mul_109_11_n_382 ^ (mul_109_11_n_925 ^ mul_109_11_n_941));
 assign mul_109_11_n_1042 = ((mul_109_11_n_988 & mul_109_11_n_922) | ((mul_109_11_n_922 & mul_109_11_n_838)
    | (mul_109_11_n_838 & mul_109_11_n_988)));
 assign mul_109_11_n_1043 = (mul_109_11_n_922 ^ (mul_109_11_n_838 ^ mul_109_11_n_988));
 assign mul_109_11_n_1040 = ((mul_109_11_n_981 & mul_109_11_n_494) | ((mul_109_11_n_494 & mul_109_11_n_910)
    | (mul_109_11_n_910 & mul_109_11_n_981)));
 assign mul_109_11_n_1041 = (mul_109_11_n_494 ^ (mul_109_11_n_910 ^ mul_109_11_n_981));
 assign mul_109_11_n_1038 = ((mul_109_11_n_915 & mul_109_11_n_507) | ((mul_109_11_n_507 & mul_109_11_n_957)
    | (mul_109_11_n_957 & mul_109_11_n_915)));
 assign mul_109_11_n_1039 = (mul_109_11_n_507 ^ (mul_109_11_n_957 ^ mul_109_11_n_915));
 assign mul_109_11_n_1036 = ((mul_109_11_n_977 & mul_109_11_n_667) | ((mul_109_11_n_667 & mul_109_11_n_859)
    | (mul_109_11_n_859 & mul_109_11_n_977)));
 assign mul_109_11_n_1037 = (mul_109_11_n_667 ^ (mul_109_11_n_859 ^ mul_109_11_n_977));
 assign mul_109_11_n_1059 = ~(mul_109_11_n_996 & mul_109_11_n_1031);
 assign mul_109_11_n_1058 = ~(mul_109_11_n_1032 & mul_109_11_n_881);
 assign {out1[7]} = ~(mul_109_11_n_1001 ^ mul_109_11_n_973);
 assign mul_109_11_n_1035 = ~(mul_109_11_n_1032 | mul_109_11_n_881);
 assign mul_109_11_n_1034 = ~(mul_109_11_n_996 | mul_109_11_n_1031);
 assign mul_109_11_n_1028 = ((mul_109_11_n_931 & mul_109_11_n_508) | ((mul_109_11_n_508 & mul_109_11_n_945)
    | (mul_109_11_n_945 & mul_109_11_n_931)));
 assign mul_109_11_n_1029 = (mul_109_11_n_508 ^ (mul_109_11_n_945 ^ mul_109_11_n_931));
 assign mul_109_11_n_1026 = ((mul_109_11_n_832 & mul_109_11_n_655) | ((mul_109_11_n_655 & mul_109_11_n_953)
    | (mul_109_11_n_953 & mul_109_11_n_832)));
 assign mul_109_11_n_1027 = (mul_109_11_n_655 ^ (mul_109_11_n_953 ^ mul_109_11_n_832));
 assign mul_109_11_n_1024 = ((mul_109_11_n_933 & mul_109_11_n_626) | ((mul_109_11_n_626 & mul_109_11_n_916)
    | (mul_109_11_n_916 & mul_109_11_n_933)));
 assign mul_109_11_n_1025 = (mul_109_11_n_626 ^ (mul_109_11_n_916 ^ mul_109_11_n_933));
 assign mul_109_11_n_1031 = ((mul_109_11_n_965 & mul_109_11_n_376) | ((mul_109_11_n_376 & mul_109_11_n_862)
    | (mul_109_11_n_862 & mul_109_11_n_965)));
 assign mul_109_11_n_1032 = (mul_109_11_n_376 ^ (mul_109_11_n_862 ^ mul_109_11_n_965));
 assign mul_109_11_n_1022 = ((mul_109_11_n_897 & mul_109_11_n_658) | ((mul_109_11_n_658 & mul_109_11_n_920)
    | (mul_109_11_n_920 & mul_109_11_n_897)));
 assign mul_109_11_n_1023 = (mul_109_11_n_658 ^ (mul_109_11_n_920 ^ mul_109_11_n_897));
 assign mul_109_11_n_1020 = ((mul_109_11_n_831 & mul_109_11_n_502) | ((mul_109_11_n_502 & mul_109_11_n_908)
    | (mul_109_11_n_908 & mul_109_11_n_831)));
 assign mul_109_11_n_1021 = (mul_109_11_n_502 ^ (mul_109_11_n_908 ^ mul_109_11_n_831));
 assign mul_109_11_n_1018 = ((mul_109_11_n_921 & mul_109_11_n_907) | ((mul_109_11_n_907 & mul_109_11_n_736)
    | (mul_109_11_n_736 & mul_109_11_n_921)));
 assign mul_109_11_n_1019 = (mul_109_11_n_907 ^ (mul_109_11_n_736 ^ mul_109_11_n_921));
 assign mul_109_11_n_1017 = ~(mul_109_11_n_998 | ~mul_109_11_n_1012);
 assign mul_109_11_n_1030 = ~(mul_109_11_n_999 | mul_109_11_n_998);
 assign mul_109_11_n_1016 = ~(mul_109_11_n_992 & (mul_109_11_n_991 | mul_109_11_n_885));
 assign mul_109_11_n_1015 = ~(mul_109_11_n_1013 & ~mul_109_11_n_999);
 assign mul_109_11_n_1014 = ~(mul_109_11_n_985 ^ mul_109_11_n_955);
 assign mul_109_11_n_1010 = ((mul_109_11_n_909 & mul_109_11_n_377) | ((mul_109_11_n_377 & mul_109_11_n_896)
    | (mul_109_11_n_896 & mul_109_11_n_909)));
 assign mul_109_11_n_1011 = (mul_109_11_n_377 ^ (mul_109_11_n_896 ^ mul_109_11_n_909));
 assign mul_109_11_n_1008 = ((mul_109_11_n_914 & mul_109_11_n_659) | ((mul_109_11_n_659 & mul_109_11_n_893)
    | (mul_109_11_n_893 & mul_109_11_n_914)));
 assign mul_109_11_n_1009 = (mul_109_11_n_659 ^ (mul_109_11_n_893 ^ mul_109_11_n_914));
 assign mul_109_11_n_1006 = ((mul_109_11_n_913 & mul_109_11_n_380) | ((mul_109_11_n_380 & mul_109_11_n_485)
    | (mul_109_11_n_485 & mul_109_11_n_913)));
 assign mul_109_11_n_1007 = (mul_109_11_n_380 ^ (mul_109_11_n_485 ^ mul_109_11_n_913));
 assign mul_109_11_n_1004 = ((mul_109_11_n_912 & mul_109_11_n_723) | ((mul_109_11_n_723 & mul_109_11_n_821)
    | (mul_109_11_n_821 & mul_109_11_n_912)));
 assign mul_109_11_n_1005 = (mul_109_11_n_723 ^ (mul_109_11_n_821 ^ mul_109_11_n_912));
 assign mul_109_11_n_1002 = ((mul_109_11_n_904 & mul_109_11_n_648) | ((mul_109_11_n_648 & mul_109_11_n_628)
    | (mul_109_11_n_628 & mul_109_11_n_904)));
 assign mul_109_11_n_1003 = (mul_109_11_n_648 ^ (mul_109_11_n_628 ^ mul_109_11_n_904));
 assign mul_109_11_n_1001 = ~(mul_109_11_n_992 & ~mul_109_11_n_991);
 assign mul_109_11_n_1013 = ~(mul_109_11_n_994 & mul_109_11_n_971);
 assign mul_109_11_n_1012 = ~(mul_109_11_n_972 & mul_109_11_n_995);
 assign mul_109_11_n_1000 = ~(mul_109_11_n_991 | mul_109_11_n_899);
 assign mul_109_11_n_997 = ~(mul_109_11_n_956 ^ mul_109_11_n_676);
 assign mul_109_11_n_999 = ~(mul_109_11_n_994 | mul_109_11_n_971);
 assign mul_109_11_n_998 = ~(mul_109_11_n_972 | mul_109_11_n_995);
 assign mul_109_11_n_989 = ((mul_109_11_n_894 & mul_109_11_n_665) | ((mul_109_11_n_665 & mul_109_11_n_778)
    | (mul_109_11_n_778 & mul_109_11_n_894)));
 assign mul_109_11_n_990 = (mul_109_11_n_665 ^ (mul_109_11_n_778 ^ mul_109_11_n_894));
 assign mul_109_11_n_995 = ((mul_109_11_n_868 & mul_109_11_n_864) | ((mul_109_11_n_864 & mul_109_11_n_810)
    | (mul_109_11_n_810 & mul_109_11_n_868)));
 assign mul_109_11_n_996 = (mul_109_11_n_864 ^ (mul_109_11_n_810 ^ mul_109_11_n_868));
 assign mul_109_11_n_993 = ((mul_109_11_n_929 & mul_109_11_n_865) | ((mul_109_11_n_865 & mul_109_11_n_725)
    | (mul_109_11_n_725 & mul_109_11_n_929)));
 assign mul_109_11_n_994 = (mul_109_11_n_865 ^ (mul_109_11_n_725 ^ mul_109_11_n_929));
 assign mul_109_11_n_987 = ((mul_109_11_n_926 & mul_109_11_n_640) | ((mul_109_11_n_640 & mul_109_11_n_841)
    | (mul_109_11_n_841 & mul_109_11_n_926)));
 assign mul_109_11_n_988 = (mul_109_11_n_640 ^ (mul_109_11_n_841 ^ mul_109_11_n_926));
 assign mul_109_11_n_985 = ((mul_109_11_n_836 & mul_109_11_n_660) | ((mul_109_11_n_660 & mul_109_11_n_890)
    | (mul_109_11_n_890 & mul_109_11_n_836)));
 assign mul_109_11_n_986 = (mul_109_11_n_660 ^ (mul_109_11_n_890 ^ mul_109_11_n_836));
 assign mul_109_11_n_983 = ((mul_109_11_n_927 & mul_109_11_n_649) | ((mul_109_11_n_649 & mul_109_11_n_842)
    | (mul_109_11_n_842 & mul_109_11_n_927)));
 assign mul_109_11_n_984 = (mul_109_11_n_649 ^ (mul_109_11_n_842 ^ mul_109_11_n_927));
 assign mul_109_11_n_981 = ((mul_109_11_n_854 & mul_109_11_n_379) | ((mul_109_11_n_379 & mul_109_11_n_856)
    | (mul_109_11_n_856 & mul_109_11_n_854)));
 assign mul_109_11_n_982 = (mul_109_11_n_379 ^ (mul_109_11_n_856 ^ mul_109_11_n_854));
 assign mul_109_11_n_979 = ((mul_109_11_n_889 & mul_109_11_n_506) | ((mul_109_11_n_506 & mul_109_11_n_654)
    | (mul_109_11_n_654 & mul_109_11_n_889)));
 assign mul_109_11_n_980 = (mul_109_11_n_506 ^ (mul_109_11_n_654 ^ mul_109_11_n_889));
 assign mul_109_11_n_977 = ((mul_109_11_n_857 & mul_109_11_n_671) | ((mul_109_11_n_671 & mul_109_11_n_852)
    | (mul_109_11_n_852 & mul_109_11_n_857)));
 assign mul_109_11_n_978 = (mul_109_11_n_671 ^ (mul_109_11_n_852 ^ mul_109_11_n_857));
 assign mul_109_11_n_975 = ((mul_109_11_n_887 & mul_109_11_n_394) | ((mul_109_11_n_394 & mul_109_11_n_782)
    | (mul_109_11_n_782 & mul_109_11_n_887)));
 assign mul_109_11_n_976 = (mul_109_11_n_394 ^ (mul_109_11_n_782 ^ mul_109_11_n_887));
 assign mul_109_11_n_992 = ~(mul_109_11_n_970 & mul_109_11_n_877);
 assign mul_109_11_n_991 = ~(mul_109_11_n_970 | mul_109_11_n_877);
 assign {out1[6]} = ~(mul_109_11_n_903 ^ mul_109_11_n_938);
 assign mul_109_11_n_973 = ~(mul_109_11_n_885 & (mul_109_11_n_938 | mul_109_11_n_899));
 assign mul_109_11_n_968 = ((mul_109_11_n_875 & mul_109_11_n_630) | ((mul_109_11_n_630 & mul_109_11_n_499)
    | (mul_109_11_n_499 & mul_109_11_n_875)));
 assign mul_109_11_n_969 = (mul_109_11_n_630 ^ (mul_109_11_n_499 ^ mul_109_11_n_875));
 assign mul_109_11_n_966 = ((mul_109_11_n_873 & mul_109_11_n_396) | ((mul_109_11_n_396 & mul_109_11_n_848)
    | (mul_109_11_n_848 & mul_109_11_n_873)));
 assign mul_109_11_n_967 = (mul_109_11_n_396 ^ (mul_109_11_n_848 ^ mul_109_11_n_873));
 assign mul_109_11_n_971 = ((mul_109_11_n_867 & mul_109_11_n_866) | ((mul_109_11_n_866 & mul_109_11_n_823)
    | (mul_109_11_n_823 & mul_109_11_n_867)));
 assign mul_109_11_n_972 = (mul_109_11_n_866 ^ (mul_109_11_n_823 ^ mul_109_11_n_867));
 assign mul_109_11_n_965 = ((mul_109_11_n_863 & mul_109_11_n_585) | ((mul_109_11_n_585 & mul_109_11_n_687)
    | (mul_109_11_n_687 & mul_109_11_n_863)));
 assign mul_109_11_n_970 = (mul_109_11_n_585 ^ (mul_109_11_n_687 ^ mul_109_11_n_863));
 assign mul_109_11_n_963 = ((mul_109_11_n_892 & mul_109_11_n_498) | ((mul_109_11_n_498 & mul_109_11_n_847)
    | (mul_109_11_n_847 & mul_109_11_n_892)));
 assign mul_109_11_n_964 = (mul_109_11_n_498 ^ (mul_109_11_n_847 ^ mul_109_11_n_892));
 assign mul_109_11_n_961 = ((mul_109_11_n_872 & mul_109_11_n_596) | ((mul_109_11_n_596 & mul_109_11_n_869)
    | (mul_109_11_n_869 & mul_109_11_n_872)));
 assign mul_109_11_n_962 = (mul_109_11_n_596 ^ (mul_109_11_n_869 ^ mul_109_11_n_872));
 assign mul_109_11_n_959 = ((mul_109_11_n_874 & mul_109_11_n_553) | ((mul_109_11_n_553 & mul_109_11_n_656)
    | (mul_109_11_n_656 & mul_109_11_n_874)));
 assign mul_109_11_n_960 = (mul_109_11_n_553 ^ (mul_109_11_n_656 ^ mul_109_11_n_874));
 assign mul_109_11_n_957 = ((mul_109_11_n_850 & mul_109_11_n_500) | ((mul_109_11_n_500 & mul_109_11_n_751)
    | (mul_109_11_n_751 & mul_109_11_n_850)));
 assign mul_109_11_n_958 = (mul_109_11_n_500 ^ (mul_109_11_n_751 ^ mul_109_11_n_850));
 assign mul_109_11_n_956 = ~(mul_109_11_n_678 ^ mul_109_11_n_924);
 assign mul_109_11_n_955 = ~(mul_109_11_n_793 ^ mul_109_11_n_919);
 assign mul_109_11_n_953 = ((mul_109_11_n_827 & mul_109_11_n_486) | ((mul_109_11_n_486 & mul_109_11_n_851)
    | (mul_109_11_n_851 & mul_109_11_n_827)));
 assign mul_109_11_n_954 = (mul_109_11_n_486 ^ (mul_109_11_n_851 ^ mul_109_11_n_827));
 assign mul_109_11_n_951 = ((mul_109_11_n_845 & mul_109_11_n_565) | ((mul_109_11_n_565 & mul_109_11_n_795)
    | (mul_109_11_n_795 & mul_109_11_n_845)));
 assign mul_109_11_n_952 = (mul_109_11_n_565 ^ (mul_109_11_n_795 ^ mul_109_11_n_845));
 assign mul_109_11_n_949 = ((mul_109_11_n_895 & mul_109_11_n_400) | ((mul_109_11_n_400 & mul_109_11_n_724)
    | (mul_109_11_n_724 & mul_109_11_n_895)));
 assign mul_109_11_n_950 = (mul_109_11_n_400 ^ (mul_109_11_n_724 ^ mul_109_11_n_895));
 assign mul_109_11_n_947 = ((mul_109_11_n_891 & mul_109_11_n_662) | ((mul_109_11_n_662 & mul_109_11_n_653)
    | (mul_109_11_n_653 & mul_109_11_n_891)));
 assign mul_109_11_n_948 = (mul_109_11_n_662 ^ (mul_109_11_n_653 ^ mul_109_11_n_891));
 assign mul_109_11_n_945 = ((mul_109_11_n_843 & mul_109_11_n_501) | ((mul_109_11_n_501 & mul_109_11_n_717)
    | (mul_109_11_n_717 & mul_109_11_n_843)));
 assign mul_109_11_n_946 = (mul_109_11_n_501 ^ (mul_109_11_n_717 ^ mul_109_11_n_843));
 assign mul_109_11_n_943 = ((mul_109_11_n_886 & mul_109_11_n_766) | ((mul_109_11_n_766 & mul_109_11_n_743)
    | (mul_109_11_n_743 & mul_109_11_n_886)));
 assign mul_109_11_n_944 = (mul_109_11_n_766 ^ (mul_109_11_n_743 ^ mul_109_11_n_886));
 assign mul_109_11_n_941 = ((mul_109_11_n_888 & mul_109_11_n_497) | ((mul_109_11_n_497 & mul_109_11_n_819)
    | (mul_109_11_n_819 & mul_109_11_n_888)));
 assign mul_109_11_n_942 = (mul_109_11_n_497 ^ (mul_109_11_n_819 ^ mul_109_11_n_888));
 assign mul_109_11_n_939 = ((mul_109_11_n_839 & mul_109_11_n_495) | ((mul_109_11_n_495 & mul_109_11_n_735)
    | (mul_109_11_n_735 & mul_109_11_n_839)));
 assign mul_109_11_n_940 = (mul_109_11_n_495 ^ (mul_109_11_n_735 ^ mul_109_11_n_839));
 assign mul_109_11_n_938 = ~(mul_109_11_n_936 | mul_109_11_n_902);
 assign {out1[5]} = ~(mul_109_11_n_901 ^ mul_109_11_n_849);
 assign mul_109_11_n_934 = ((mul_109_11_n_853 & mul_109_11_n_401) | ((mul_109_11_n_401 & mul_109_11_n_627)
    | (mul_109_11_n_627 & mul_109_11_n_853)));
 assign mul_109_11_n_935 = (mul_109_11_n_401 ^ (mul_109_11_n_627 ^ mul_109_11_n_853));
 assign mul_109_11_n_932 = ((mul_109_11_n_758 & mul_109_11_n_666) | ((mul_109_11_n_666 & mul_109_11_n_798)
    | (mul_109_11_n_798 & mul_109_11_n_758)));
 assign mul_109_11_n_933 = (mul_109_11_n_666 ^ (mul_109_11_n_798 ^ mul_109_11_n_758));
 assign mul_109_11_n_930 = ((mul_109_11_n_785 & mul_109_11_n_840) | ((mul_109_11_n_840 & mul_109_11_n_756)
    | (mul_109_11_n_756 & mul_109_11_n_785)));
 assign mul_109_11_n_931 = (mul_109_11_n_840 ^ (mul_109_11_n_756 ^ mul_109_11_n_785));
 assign mul_109_11_n_928 = ((mul_109_11_n_822 & mul_109_11_n_444) | ((mul_109_11_n_444 & mul_109_11_n_825)
    | (mul_109_11_n_825 & mul_109_11_n_822)));
 assign mul_109_11_n_929 = (mul_109_11_n_444 ^ (mul_109_11_n_825 ^ mul_109_11_n_822));
 assign mul_109_11_n_926 = ((mul_109_11_n_803 & mul_109_11_n_582) | ((mul_109_11_n_582 & mul_109_11_n_805)
    | (mul_109_11_n_805 & mul_109_11_n_803)));
 assign mul_109_11_n_927 = (mul_109_11_n_582 ^ (mul_109_11_n_805 ^ mul_109_11_n_803));
 assign mul_109_11_n_924 = ((mul_109_11_n_762 & mul_109_11_n_503) | ((mul_109_11_n_503 & mul_109_11_n_818)
    | (mul_109_11_n_818 & mul_109_11_n_762)));
 assign mul_109_11_n_925 = (mul_109_11_n_503 ^ (mul_109_11_n_818 ^ mul_109_11_n_762));
 assign mul_109_11_n_922 = ((mul_109_11_n_858 & mul_109_11_n_551) | ((mul_109_11_n_551 & mul_109_11_n_637)
    | (mul_109_11_n_637 & mul_109_11_n_858)));
 assign mul_109_11_n_923 = (mul_109_11_n_551 ^ (mul_109_11_n_637 ^ mul_109_11_n_858));
 assign mul_109_11_n_920 = ((mul_109_11_n_820 & mul_109_11_n_641) | ((mul_109_11_n_641 & mul_109_11_n_789)
    | (mul_109_11_n_789 & mul_109_11_n_820)));
 assign mul_109_11_n_921 = (mul_109_11_n_641 ^ (mul_109_11_n_789 ^ mul_109_11_n_820));
 assign mul_109_11_n_936 = ~(mul_109_11_n_900 & (mul_109_11_n_898 | mul_109_11_n_816));
 assign mul_109_11_n_919 = ~(mul_109_11_n_860 ^ mul_109_11_n_883);
 assign mul_109_11_n_918 = ~(mul_109_11_n_543 ^ mul_109_11_n_882);
 assign mul_109_11_n_916 = ((mul_109_11_n_799 & mul_109_11_n_555) | ((mul_109_11_n_555 & mul_109_11_n_398)
    | (mul_109_11_n_398 & mul_109_11_n_799)));
 assign mul_109_11_n_917 = (mul_109_11_n_555 ^ (mul_109_11_n_398 ^ mul_109_11_n_799));
 assign mul_109_11_n_914 = ((mul_109_11_n_844 & mul_109_11_n_492) | ((mul_109_11_n_492 & mul_109_11_n_750)
    | (mul_109_11_n_750 & mul_109_11_n_844)));
 assign mul_109_11_n_915 = (mul_109_11_n_492 ^ (mul_109_11_n_750 ^ mul_109_11_n_844));
 assign mul_109_11_n_912 = ((mul_109_11_n_802 & mul_109_11_n_528) | ((mul_109_11_n_528 & mul_109_11_n_772)
    | (mul_109_11_n_772 & mul_109_11_n_802)));
 assign mul_109_11_n_913 = (mul_109_11_n_528 ^ (mul_109_11_n_772 ^ mul_109_11_n_802));
 assign mul_109_11_n_910 = ((mul_109_11_n_806 & mul_109_11_n_635) | ((mul_109_11_n_635 & mul_109_11_n_618)
    | (mul_109_11_n_618 & mul_109_11_n_806)));
 assign mul_109_11_n_911 = (mul_109_11_n_635 ^ (mul_109_11_n_618 ^ mul_109_11_n_806));
 assign mul_109_11_n_908 = ((mul_109_11_n_826 & mul_109_11_n_780) | ((mul_109_11_n_780 & mul_109_11_n_749)
    | (mul_109_11_n_749 & mul_109_11_n_826)));
 assign mul_109_11_n_909 = (mul_109_11_n_780 ^ (mul_109_11_n_749 ^ mul_109_11_n_826));
 assign mul_109_11_n_906 = ((mul_109_11_n_811 & mul_109_11_n_397) | ((mul_109_11_n_397 & mul_109_11_n_484)
    | (mul_109_11_n_484 & mul_109_11_n_811)));
 assign mul_109_11_n_907 = (mul_109_11_n_397 ^ (mul_109_11_n_484 ^ mul_109_11_n_811));
 assign mul_109_11_n_904 = ((mul_109_11_n_794 & mul_109_11_n_580) | ((mul_109_11_n_580 & mul_109_11_n_739)
    | (mul_109_11_n_739 & mul_109_11_n_794)));
 assign mul_109_11_n_905 = (mul_109_11_n_580 ^ (mul_109_11_n_739 ^ mul_109_11_n_794));
 assign mul_109_11_n_903 = ~(mul_109_11_n_899 | ~mul_109_11_n_885);
 assign mul_109_11_n_901 = ~(mul_109_11_n_900 & ~mul_109_11_n_898);
 assign mul_109_11_n_902 = ~(mul_109_11_n_898 | mul_109_11_n_829);
 assign mul_109_11_n_896 = ((mul_109_11_n_788 & mul_109_11_n_644) | ((mul_109_11_n_644 & mul_109_11_n_781)
    | (mul_109_11_n_781 & mul_109_11_n_788)));
 assign mul_109_11_n_897 = (mul_109_11_n_644 ^ (mul_109_11_n_781 ^ mul_109_11_n_788));
 assign mul_109_11_n_894 = ((mul_109_11_n_824 & mul_109_11_n_445) | ((mul_109_11_n_445 & mul_109_11_n_702)
    | (mul_109_11_n_702 & mul_109_11_n_824)));
 assign mul_109_11_n_895 = (mul_109_11_n_445 ^ (mul_109_11_n_702 ^ mul_109_11_n_824));
 assign mul_109_11_n_892 = ((mul_109_11_n_786 & mul_109_11_n_487) | ((mul_109_11_n_487 & mul_109_11_n_764)
    | (mul_109_11_n_764 & mul_109_11_n_786)));
 assign mul_109_11_n_893 = (mul_109_11_n_487 ^ (mul_109_11_n_764 ^ mul_109_11_n_786));
 assign mul_109_11_n_890 = ((mul_109_11_n_790 & mul_109_11_n_483) | ((mul_109_11_n_483 & mul_109_11_n_734)
    | (mul_109_11_n_734 & mul_109_11_n_790)));
 assign mul_109_11_n_891 = (mul_109_11_n_483 ^ (mul_109_11_n_734 ^ mul_109_11_n_790));
 assign mul_109_11_n_888 = ((mul_109_11_n_791 & mul_109_11_n_490) | ((mul_109_11_n_490 & mul_109_11_n_784)
    | (mul_109_11_n_784 & mul_109_11_n_791)));
 assign mul_109_11_n_889 = (mul_109_11_n_490 ^ (mul_109_11_n_784 ^ mul_109_11_n_791));
 assign mul_109_11_n_886 = ((mul_109_11_n_721 & mul_109_11_n_651) | ((mul_109_11_n_651 & mul_109_11_n_755)
    | (mul_109_11_n_755 & mul_109_11_n_721)));
 assign mul_109_11_n_887 = (mul_109_11_n_651 ^ (mul_109_11_n_755 ^ mul_109_11_n_721));
 assign mul_109_11_n_900 = ~(mul_109_11_n_880 & mul_109_11_n_615);
 assign mul_109_11_n_899 = ~(mul_109_11_n_878 | mul_109_11_n_879);
 assign mul_109_11_n_898 = ~(mul_109_11_n_880 | mul_109_11_n_615);
 assign {out1[4]} = ~(mul_109_11_n_830 ^ mul_109_11_n_814);
 assign mul_109_11_n_883 = ~(mul_109_11_n_779 ^ mul_109_11_n_835);
 assign mul_109_11_n_882 = ~(mul_109_11_n_675 ^ mul_109_11_n_828);
 assign mul_109_11_n_885 = ~(mul_109_11_n_878 & mul_109_11_n_879);
 assign mul_109_11_n_875 = ((mul_109_11_n_797 & mul_109_11_n_634) | ((mul_109_11_n_634 & mul_109_11_n_722)
    | (mul_109_11_n_722 & mul_109_11_n_797)));
 assign mul_109_11_n_876 = (mul_109_11_n_634 ^ (mul_109_11_n_722 ^ mul_109_11_n_797));
 assign mul_109_11_n_873 = ((mul_109_11_n_787 & mul_109_11_n_652) | ((mul_109_11_n_652 & mul_109_11_n_731)
    | (mul_109_11_n_731 & mul_109_11_n_787)));
 assign mul_109_11_n_874 = (mul_109_11_n_652 ^ (mul_109_11_n_731 ^ mul_109_11_n_787));
 assign mul_109_11_n_871 = ((mul_109_11_n_775 & mul_109_11_n_436) | ((mul_109_11_n_436 & mul_109_11_n_496)
    | (mul_109_11_n_496 & mul_109_11_n_775)));
 assign mul_109_11_n_872 = (mul_109_11_n_436 ^ (mul_109_11_n_496 ^ mul_109_11_n_775));
 assign mul_109_11_n_869 = ((mul_109_11_n_776 & mul_109_11_n_437) | ((mul_109_11_n_437 & mul_109_11_n_482)
    | (mul_109_11_n_482 & mul_109_11_n_776)));
 assign mul_109_11_n_870 = (mul_109_11_n_437 ^ (mul_109_11_n_482 ^ mul_109_11_n_776));
 assign mul_109_11_n_867 = ((mul_109_11_n_773 & mul_109_11_n_454) | ((mul_109_11_n_454 & mul_109_11_n_395)
    | (mul_109_11_n_395 & mul_109_11_n_773)));
 assign mul_109_11_n_868 = (mul_109_11_n_454 ^ (mul_109_11_n_395 ^ mul_109_11_n_773));
 assign mul_109_11_n_865 = ((mul_109_11_n_809 & mul_109_11_n_378) | ((mul_109_11_n_378 & mul_109_11_n_443)
    | (mul_109_11_n_443 & mul_109_11_n_809)));
 assign mul_109_11_n_866 = (mul_109_11_n_378 ^ (mul_109_11_n_443 ^ mul_109_11_n_809));
 assign mul_109_11_n_864 = ((mul_109_11_n_774 & mul_109_11_n_584) | ((mul_109_11_n_584 & mul_109_11_n_518)
    | (mul_109_11_n_518 & mul_109_11_n_774)));
 assign mul_109_11_n_881 = (mul_109_11_n_584 ^ (mul_109_11_n_518 ^ mul_109_11_n_774));
 assign mul_109_11_n_862 = ((mul_109_11_n_807 & mul_109_11_n_664) | ((mul_109_11_n_664 & mul_109_11_n_561)
    | (mul_109_11_n_561 & mul_109_11_n_807)));
 assign mul_109_11_n_863 = (mul_109_11_n_664 ^ (mul_109_11_n_561 ^ mul_109_11_n_807));
 assign mul_109_11_n_879 = ((mul_109_11_n_813 & mul_109_11_n_701) | ((mul_109_11_n_701 & mul_109_11_n_415)
    | (mul_109_11_n_415 & mul_109_11_n_813)));
 assign mul_109_11_n_880 = (mul_109_11_n_701 ^ (mul_109_11_n_415 ^ mul_109_11_n_813));
 assign mul_109_11_n_877 = ((mul_109_11_n_808 & mul_109_11_n_403) | ((mul_109_11_n_403 & mul_109_11_n_556)
    | (mul_109_11_n_556 & mul_109_11_n_808)));
 assign mul_109_11_n_878 = (mul_109_11_n_403 ^ (mul_109_11_n_556 ^ mul_109_11_n_808));
 assign mul_109_11_n_860 = ((mul_109_11_n_765 & mul_109_11_n_491) | ((mul_109_11_n_491 & mul_109_11_n_770)
    | (mul_109_11_n_770 & mul_109_11_n_765)));
 assign mul_109_11_n_861 = (mul_109_11_n_491 ^ (mul_109_11_n_770 ^ mul_109_11_n_765));
 assign mul_109_11_n_858 = ((mul_109_11_n_800 & mul_109_11_n_526) | ((mul_109_11_n_526 & mul_109_11_n_747)
    | (mul_109_11_n_747 & mul_109_11_n_800)));
 assign mul_109_11_n_859 = (mul_109_11_n_526 ^ (mul_109_11_n_747 ^ mul_109_11_n_800));
 assign mul_109_11_n_856 = ((mul_109_11_n_759 & mul_109_11_n_524) | ((mul_109_11_n_524 & mul_109_11_n_416)
    | (mul_109_11_n_416 & mul_109_11_n_759)));
 assign mul_109_11_n_857 = (mul_109_11_n_524 ^ (mul_109_11_n_416 ^ mul_109_11_n_759));
 assign mul_109_11_n_854 = ((mul_109_11_n_801 & mul_109_11_n_617) | ((mul_109_11_n_617 & mul_109_11_n_738)
    | (mul_109_11_n_738 & mul_109_11_n_801)));
 assign mul_109_11_n_855 = (mul_109_11_n_617 ^ (mul_109_11_n_738 ^ mul_109_11_n_801));
 assign mul_109_11_n_852 = ((mul_109_11_n_760 & mul_109_11_n_517) | ((mul_109_11_n_517 & mul_109_11_n_757)
    | (mul_109_11_n_757 & mul_109_11_n_760)));
 assign mul_109_11_n_853 = (mul_109_11_n_517 ^ (mul_109_11_n_757 ^ mul_109_11_n_760));
 assign mul_109_11_n_850 = ((mul_109_11_n_796 & mul_109_11_n_632) | ((mul_109_11_n_632 & mul_109_11_n_512)
    | (mul_109_11_n_512 & mul_109_11_n_796)));
 assign mul_109_11_n_851 = (mul_109_11_n_632 ^ (mul_109_11_n_512 ^ mul_109_11_n_796));
 assign mul_109_11_n_849 = ~(mul_109_11_n_829 & mul_109_11_n_816);
 assign mul_109_11_n_847 = ((mul_109_11_n_727 & mul_109_11_n_643) | ((mul_109_11_n_643 & mul_109_11_n_730)
    | (mul_109_11_n_730 & mul_109_11_n_727)));
 assign mul_109_11_n_848 = (mul_109_11_n_643 ^ (mul_109_11_n_730 ^ mul_109_11_n_727));
 assign mul_109_11_n_845 = ((mul_109_11_n_753 & mul_109_11_n_431) | ((mul_109_11_n_431 & mul_109_11_n_777)
    | (mul_109_11_n_777 & mul_109_11_n_753)));
 assign mul_109_11_n_846 = (mul_109_11_n_431 ^ (mul_109_11_n_777 ^ mul_109_11_n_753));
 assign mul_109_11_n_843 = ((mul_109_11_n_748 & mul_109_11_n_516) | ((mul_109_11_n_516 & mul_109_11_n_740)
    | (mul_109_11_n_740 & mul_109_11_n_748)));
 assign mul_109_11_n_844 = (mul_109_11_n_516 ^ (mul_109_11_n_740 ^ mul_109_11_n_748));
 assign mul_109_11_n_841 = ((mul_109_11_n_746 & mul_109_11_n_529) | ((mul_109_11_n_529 & mul_109_11_n_427)
    | (mul_109_11_n_427 & mul_109_11_n_746)));
 assign mul_109_11_n_842 = (mul_109_11_n_529 ^ (mul_109_11_n_427 ^ mul_109_11_n_746));
 assign mul_109_11_n_839 = ((mul_109_11_n_763 & mul_109_11_n_531) | ((mul_109_11_n_531 & mul_109_11_n_726)
    | (mul_109_11_n_726 & mul_109_11_n_763)));
 assign mul_109_11_n_840 = (mul_109_11_n_531 ^ (mul_109_11_n_726 ^ mul_109_11_n_763));
 assign mul_109_11_n_837 = ((mul_109_11_n_729 & mul_109_11_n_638) | ((mul_109_11_n_638 & mul_109_11_n_549)
    | (mul_109_11_n_549 & mul_109_11_n_729)));
 assign mul_109_11_n_838 = (mul_109_11_n_638 ^ (mul_109_11_n_549 ^ mul_109_11_n_729));
 assign mul_109_11_n_835 = ((mul_109_11_n_745 & mul_109_11_n_650) | ((mul_109_11_n_650 & mul_109_11_n_742)
    | (mul_109_11_n_742 & mul_109_11_n_745)));
 assign mul_109_11_n_836 = (mul_109_11_n_650 ^ (mul_109_11_n_742 ^ mul_109_11_n_745));
 assign mul_109_11_n_833 = ((mul_109_11_n_783 & mul_109_11_n_661) | ((mul_109_11_n_661 & mul_109_11_n_657)
    | (mul_109_11_n_657 & mul_109_11_n_783)));
 assign mul_109_11_n_834 = (mul_109_11_n_661 ^ (mul_109_11_n_657 ^ mul_109_11_n_783));
 assign mul_109_11_n_831 = ((mul_109_11_n_741 & mul_109_11_n_489) | ((mul_109_11_n_489 & mul_109_11_n_647)
    | (mul_109_11_n_647 & mul_109_11_n_741)));
 assign mul_109_11_n_832 = (mul_109_11_n_489 ^ (mul_109_11_n_647 ^ mul_109_11_n_741));
 assign mul_109_11_n_830 = ~(mul_109_11_n_816 & ~mul_109_11_n_817);
 assign mul_109_11_n_829 = ~(mul_109_11_n_814 & ~mul_109_11_n_817);
 assign mul_109_11_n_828 = ~(mul_109_11_n_792 ^ mul_109_11_n_769);
 assign mul_109_11_n_826 = ((mul_109_11_n_718 & mul_109_11_n_432) | ((mul_109_11_n_432 & mul_109_11_n_575)
    | (mul_109_11_n_575 & mul_109_11_n_718)));
 assign mul_109_11_n_827 = (mul_109_11_n_432 ^ (mul_109_11_n_575 ^ mul_109_11_n_718));
 assign mul_109_11_n_824 = ((mul_109_11_n_767 & mul_109_11_n_589) | ((mul_109_11_n_589 & mul_109_11_n_703)
    | (mul_109_11_n_703 & mul_109_11_n_767)));
 assign mul_109_11_n_825 = (mul_109_11_n_589 ^ (mul_109_11_n_703 ^ mul_109_11_n_767));
 assign mul_109_11_n_822 = ((mul_109_11_n_768 & mul_109_11_n_586) | ((mul_109_11_n_586 & mul_109_11_n_532)
    | (mul_109_11_n_532 & mul_109_11_n_768)));
 assign mul_109_11_n_823 = (mul_109_11_n_586 ^ (mul_109_11_n_532 ^ mul_109_11_n_768));
 assign mul_109_11_n_820 = ((mul_109_11_n_771 & mul_109_11_n_579) | ((mul_109_11_n_579 & mul_109_11_n_699)
    | (mul_109_11_n_699 & mul_109_11_n_771)));
 assign mul_109_11_n_821 = (mul_109_11_n_579 ^ (mul_109_11_n_699 ^ mul_109_11_n_771));
 assign mul_109_11_n_818 = ((mul_109_11_n_720 & mul_109_11_n_645) | ((mul_109_11_n_645 & mul_109_11_n_515)
    | (mul_109_11_n_515 & mul_109_11_n_720)));
 assign mul_109_11_n_819 = (mul_109_11_n_645 ^ (mul_109_11_n_515 ^ mul_109_11_n_720));
 assign mul_109_11_n_817 = ~(mul_109_11_n_815 | mul_109_11_n_480);
 assign mul_109_11_n_816 = ~(mul_109_11_n_815 & mul_109_11_n_480);
 assign mul_109_11_n_813 = ((mul_109_11_n_694 & mul_109_11_n_399) | ((mul_109_11_n_399 & mul_109_11_n_523)
    | (mul_109_11_n_523 & mul_109_11_n_694)));
 assign mul_109_11_n_815 = (mul_109_11_n_399 ^ (mul_109_11_n_523 ^ mul_109_11_n_694));
 assign mul_109_11_n_811 = ((mul_109_11_n_728 & mul_109_11_n_623) | ((mul_109_11_n_623 & mul_109_11_n_525)
    | (mul_109_11_n_525 & mul_109_11_n_728)));
 assign mul_109_11_n_812 = (mul_109_11_n_623 ^ (mul_109_11_n_525 ^ mul_109_11_n_728));
 assign mul_109_11_n_809 = ((mul_109_11_n_707 & mul_109_11_n_587) | ((mul_109_11_n_587 & mul_109_11_n_533)
    | (mul_109_11_n_533 & mul_109_11_n_707)));
 assign mul_109_11_n_810 = (mul_109_11_n_587 ^ (mul_109_11_n_533 ^ mul_109_11_n_707));
 assign mul_109_11_n_807 = ((mul_109_11_n_700 & mul_109_11_n_530) | ((mul_109_11_n_530 & mul_109_11_n_419)
    | (mul_109_11_n_419 & mul_109_11_n_700)));
 assign mul_109_11_n_808 = (mul_109_11_n_530 ^ (mul_109_11_n_419 ^ mul_109_11_n_700));
 assign mul_109_11_n_805 = ((mul_109_11_n_708 & mul_109_11_n_414) | ((mul_109_11_n_414 & mul_109_11_n_423)
    | (mul_109_11_n_423 & mul_109_11_n_708)));
 assign mul_109_11_n_806 = (mul_109_11_n_414 ^ (mul_109_11_n_423 ^ mul_109_11_n_708));
 assign mul_109_11_n_814 = ((mul_109_11_n_732 & mul_109_11_n_478) | ((mul_109_11_n_478 & mul_109_11_n_695)
    | (mul_109_11_n_695 & mul_109_11_n_732)));
 assign {out1[3]} = (mul_109_11_n_478 ^ (mul_109_11_n_695 ^ mul_109_11_n_732));
 assign mul_109_11_n_802 = ((mul_109_11_n_713 & mul_109_11_n_481) | ((mul_109_11_n_481 & mul_109_11_n_578)
    | (mul_109_11_n_578 & mul_109_11_n_713)));
 assign mul_109_11_n_803 = (mul_109_11_n_481 ^ (mul_109_11_n_578 ^ mul_109_11_n_713));
 assign mul_109_11_n_800 = ((mul_109_11_n_709 & mul_109_11_n_438) | ((mul_109_11_n_438 & mul_109_11_n_576)
    | (mul_109_11_n_576 & mul_109_11_n_709)));
 assign mul_109_11_n_801 = (mul_109_11_n_438 ^ (mul_109_11_n_576 ^ mul_109_11_n_709));
 assign mul_109_11_n_798 = ((mul_109_11_n_710 & mul_109_11_n_513) | ((mul_109_11_n_513 & mul_109_11_n_430)
    | (mul_109_11_n_430 & mul_109_11_n_710)));
 assign mul_109_11_n_799 = (mul_109_11_n_513 ^ (mul_109_11_n_430 ^ mul_109_11_n_710));
 assign mul_109_11_n_796 = ((mul_109_11_n_698 & mul_109_11_n_417) | ((mul_109_11_n_417 & mul_109_11_n_567)
    | (mul_109_11_n_567 & mul_109_11_n_698)));
 assign mul_109_11_n_797 = (mul_109_11_n_417 ^ (mul_109_11_n_567 ^ mul_109_11_n_698));
 assign mul_109_11_n_794 = ((mul_109_11_n_752 & mul_109_11_n_425) | ((mul_109_11_n_425 & mul_109_11_n_514)
    | (mul_109_11_n_514 & mul_109_11_n_752)));
 assign mul_109_11_n_795 = (mul_109_11_n_425 ^ (mul_109_11_n_514 ^ mul_109_11_n_752));
 assign mul_109_11_n_793 = ~(mul_109_11_n_542 ^ mul_109_11_n_754);
 assign mul_109_11_n_792 = ~(mul_109_11_n_541 ^ mul_109_11_n_761);
 assign mul_109_11_n_790 = ((mul_109_11_n_690 & mul_109_11_n_519) | ((mul_109_11_n_519 & mul_109_11_n_588)
    | (mul_109_11_n_588 & mul_109_11_n_690)));
 assign mul_109_11_n_791 = (mul_109_11_n_519 ^ (mul_109_11_n_588 ^ mul_109_11_n_690));
 assign mul_109_11_n_788 = ((mul_109_11_n_719 & mul_109_11_n_527) | ((mul_109_11_n_527 & mul_109_11_n_594)
    | (mul_109_11_n_594 & mul_109_11_n_719)));
 assign mul_109_11_n_789 = (mul_109_11_n_527 ^ (mul_109_11_n_594 ^ mul_109_11_n_719));
 assign mul_109_11_n_786 = ((mul_109_11_n_693 & mul_109_11_n_624) | ((mul_109_11_n_624 & mul_109_11_n_571)
    | (mul_109_11_n_571 & mul_109_11_n_693)));
 assign mul_109_11_n_787 = (mul_109_11_n_624 ^ (mul_109_11_n_571 ^ mul_109_11_n_693));
 assign mul_109_11_n_784 = ((mul_109_11_n_691 & mul_109_11_n_429) | ((mul_109_11_n_429 & mul_109_11_n_636)
    | (mul_109_11_n_636 & mul_109_11_n_691)));
 assign mul_109_11_n_785 = (mul_109_11_n_429 ^ (mul_109_11_n_636 ^ mul_109_11_n_691));
 assign mul_109_11_n_782 = ((mul_109_11_n_716 & mul_109_11_n_488) | ((mul_109_11_n_488 & mul_109_11_n_646)
    | (mul_109_11_n_646 & mul_109_11_n_716)));
 assign mul_109_11_n_783 = (mul_109_11_n_488 ^ (mul_109_11_n_646 ^ mul_109_11_n_716));
 assign mul_109_11_n_780 = ((mul_109_11_n_689 & mul_109_11_n_569) | ((mul_109_11_n_569 & mul_109_11_n_595)
    | (mul_109_11_n_595 & mul_109_11_n_689)));
 assign mul_109_11_n_781 = (mul_109_11_n_569 ^ (mul_109_11_n_595 ^ mul_109_11_n_689));
 assign mul_109_11_n_779 = ~(mul_109_11_n_682 ^ mul_109_11_n_744);
 assign mul_109_11_n_777 = ((mul_109_11_n_711 & mul_109_11_n_439) | ((mul_109_11_n_439 & mul_109_11_n_428)
    | (mul_109_11_n_428 & mul_109_11_n_711)));
 assign mul_109_11_n_778 = (mul_109_11_n_439 ^ (mul_109_11_n_428 ^ mul_109_11_n_711));
 assign mul_109_11_n_775 = ((mul_109_11_n_473 & mul_109_11_n_590) | ((mul_109_11_n_590 & mul_109_11_n_566)
    | (mul_109_11_n_566 & mul_109_11_n_473)));
 assign mul_109_11_n_776 = (mul_109_11_n_590 ^ (mul_109_11_n_566 ^ mul_109_11_n_473));
 assign mul_109_11_n_773 = ((mul_109_11_n_686 & mul_109_11_n_559) | ((mul_109_11_n_559 & mul_109_11_n_421)
    | (mul_109_11_n_421 & mul_109_11_n_686)));
 assign mul_109_11_n_774 = (mul_109_11_n_559 ^ (mul_109_11_n_421 ^ mul_109_11_n_686));
 assign mul_109_11_n_771 = ((mul_109_11_n_712 & mul_109_11_n_442) | ((mul_109_11_n_442 & mul_109_11_n_581)
    | (mul_109_11_n_581 & mul_109_11_n_712)));
 assign mul_109_11_n_772 = (mul_109_11_n_442 ^ (mul_109_11_n_581 ^ mul_109_11_n_712));
 assign mul_109_11_n_769 = ((mul_109_11_n_540 & mul_109_11_n_633) | ((mul_109_11_n_633 & mul_109_11_n_554)
    | (mul_109_11_n_554 & mul_109_11_n_540)));
 assign mul_109_11_n_770 = (mul_109_11_n_633 ^ (mul_109_11_n_554 ^ mul_109_11_n_540));
 assign mul_109_11_n_767 = ((mul_109_11_n_706 & mul_109_11_n_424) | ((mul_109_11_n_424 & mul_109_11_n_564)
    | (mul_109_11_n_564 & mul_109_11_n_706)));
 assign mul_109_11_n_768 = (mul_109_11_n_424 ^ (mul_109_11_n_564 ^ mul_109_11_n_706));
 assign mul_109_11_n_765 = ((mul_109_11_n_705 & mul_109_11_n_520) | ((mul_109_11_n_520 & mul_109_11_n_558)
    | (mul_109_11_n_558 & mul_109_11_n_705)));
 assign mul_109_11_n_766 = (mul_109_11_n_520 ^ (mul_109_11_n_558 ^ mul_109_11_n_705));
 assign mul_109_11_n_763 = ((mul_109_11_n_692 & mul_109_11_n_563) | ((mul_109_11_n_563 & mul_109_11_n_591)
    | (mul_109_11_n_591 & mul_109_11_n_692)));
 assign mul_109_11_n_764 = (mul_109_11_n_563 ^ (mul_109_11_n_591 ^ mul_109_11_n_692));
 assign mul_109_11_n_761 = ((mul_109_11_n_704 & mul_109_11_n_521) | ((mul_109_11_n_521 & mul_109_11_n_663)
    | (mul_109_11_n_663 & mul_109_11_n_704)));
 assign mul_109_11_n_762 = (mul_109_11_n_521 ^ (mul_109_11_n_663 ^ mul_109_11_n_704));
 assign mul_109_11_n_759 = ((mul_109_11_n_696 & mul_109_11_n_434) | ((mul_109_11_n_434 & mul_109_11_n_557)
    | (mul_109_11_n_557 & mul_109_11_n_696)));
 assign mul_109_11_n_760 = (mul_109_11_n_434 ^ (mul_109_11_n_557 ^ mul_109_11_n_696));
 assign mul_109_11_n_757 = ((mul_109_11_n_697 & mul_109_11_n_455) | ((mul_109_11_n_455 & mul_109_11_n_452)
    | (mul_109_11_n_452 & mul_109_11_n_697)));
 assign mul_109_11_n_758 = (mul_109_11_n_455 ^ (mul_109_11_n_452 ^ mul_109_11_n_697));
 assign mul_109_11_n_755 = ((mul_109_11_n_611 & mul_109_11_n_621) | ((mul_109_11_n_621 & mul_109_11_n_577)
    | (mul_109_11_n_577 & mul_109_11_n_611)));
 assign mul_109_11_n_756 = (mul_109_11_n_621 ^ (mul_109_11_n_577 ^ mul_109_11_n_611));
 assign mul_109_11_n_754 = ~(mul_109_11_n_714 ^ mul_109_11_n_715);
 assign mul_109_11_n_752 = ((mul_109_11_n_609 & mul_109_11_n_450) | ((mul_109_11_n_450 & mul_109_11_n_570)
    | (mul_109_11_n_570 & mul_109_11_n_609)));
 assign mul_109_11_n_753 = (mul_109_11_n_450 ^ (mul_109_11_n_570 ^ mul_109_11_n_609));
 assign mul_109_11_n_750 = ((mul_109_11_n_674 & mul_109_11_n_522) | ((mul_109_11_n_522 & mul_109_11_n_435)
    | (mul_109_11_n_435 & mul_109_11_n_674)));
 assign mul_109_11_n_751 = (mul_109_11_n_522 ^ (mul_109_11_n_435 ^ mul_109_11_n_674));
 assign mul_109_11_n_748 = ((mul_109_11_n_688 & mul_109_11_n_451) | ((mul_109_11_n_451 & mul_109_11_n_449)
    | (mul_109_11_n_449 & mul_109_11_n_688)));
 assign mul_109_11_n_749 = (mul_109_11_n_451 ^ (mul_109_11_n_449 ^ mul_109_11_n_688));
 assign mul_109_11_n_746 = ((mul_109_11_n_598 & mul_109_11_n_562) | ((mul_109_11_n_562 & mul_109_11_n_440)
    | (mul_109_11_n_440 & mul_109_11_n_598)));
 assign mul_109_11_n_747 = (mul_109_11_n_562 ^ (mul_109_11_n_440 ^ mul_109_11_n_598));
 assign mul_109_11_n_744 = ((mul_109_11_n_673 & mul_109_11_n_453) | ((mul_109_11_n_453 & mul_109_11_n_413)
    | (mul_109_11_n_413 & mul_109_11_n_673)));
 assign mul_109_11_n_745 = (mul_109_11_n_453 ^ (mul_109_11_n_413 ^ mul_109_11_n_673));
 assign mul_109_11_n_742 = ((mul_109_11_n_470 & mul_109_11_n_625) | ((mul_109_11_n_625 & mul_109_11_n_583)
    | (mul_109_11_n_583 & mul_109_11_n_470)));
 assign mul_109_11_n_743 = (mul_109_11_n_625 ^ (mul_109_11_n_583 ^ mul_109_11_n_470));
 assign mul_109_11_n_740 = ((mul_109_11_n_610 & mul_109_11_n_572) | ((mul_109_11_n_572 & mul_109_11_n_616)
    | (mul_109_11_n_616 & mul_109_11_n_610)));
 assign mul_109_11_n_741 = (mul_109_11_n_572 ^ (mul_109_11_n_616 ^ mul_109_11_n_610));
 assign mul_109_11_n_738 = ((mul_109_11_n_471 & mul_109_11_n_420) | ((mul_109_11_n_420 & mul_109_11_n_574)
    | (mul_109_11_n_574 & mul_109_11_n_471)));
 assign mul_109_11_n_739 = (mul_109_11_n_420 ^ (mul_109_11_n_574 ^ mul_109_11_n_471));
 assign mul_109_11_n_736 = ((mul_109_11_n_535 & mul_109_11_n_552) | ((mul_109_11_n_552 & mul_109_11_n_642)
    | (mul_109_11_n_642 & mul_109_11_n_535)));
 assign mul_109_11_n_737 = (mul_109_11_n_552 ^ (mul_109_11_n_642 ^ mul_109_11_n_535));
 assign mul_109_11_n_734 = ((mul_109_11_n_539 & mul_109_11_n_631) | ((mul_109_11_n_631 & mul_109_11_n_573)
    | (mul_109_11_n_573 & mul_109_11_n_539)));
 assign mul_109_11_n_735 = (mul_109_11_n_631 ^ (mul_109_11_n_573 ^ mul_109_11_n_539));
 assign mul_109_11_n_732 = ((mul_109_11_n_680 & mul_109_11_n_381) | ((mul_109_11_n_381 & mul_109_11_n_544)
    | (mul_109_11_n_544 & mul_109_11_n_680)));
 assign {out1[2]} = (mul_109_11_n_381 ^ (mul_109_11_n_544 ^ mul_109_11_n_680));
 assign mul_109_11_n_730 = ((mul_109_11_n_600 & mul_109_11_n_418) | ((mul_109_11_n_418 & mul_109_11_n_568)
    | (mul_109_11_n_568 & mul_109_11_n_600)));
 assign mul_109_11_n_731 = (mul_109_11_n_418 ^ (mul_109_11_n_568 ^ mul_109_11_n_600));
 assign mul_109_11_n_728 = ((mul_109_11_n_599 & mul_109_11_n_433) | ((mul_109_11_n_433 & mul_109_11_n_446)
    | (mul_109_11_n_446 & mul_109_11_n_599)));
 assign mul_109_11_n_729 = (mul_109_11_n_433 ^ (mul_109_11_n_446 ^ mul_109_11_n_599));
 assign mul_109_11_n_726 = ((mul_109_11_n_457 & mul_109_11_n_592) | ((mul_109_11_n_592 & mul_109_11_n_448)
    | (mul_109_11_n_448 & mul_109_11_n_457)));
 assign mul_109_11_n_727 = (mul_109_11_n_592 ^ (mul_109_11_n_448 ^ mul_109_11_n_457));
 assign mul_109_11_n_724 = ((mul_109_11_n_466 & mul_109_11_n_550) | ((mul_109_11_n_550 & mul_109_11_n_493)
    | (mul_109_11_n_493 & mul_109_11_n_466)));
 assign mul_109_11_n_725 = (mul_109_11_n_550 ^ (mul_109_11_n_493 ^ mul_109_11_n_466));
 assign mul_109_11_n_722 = ((mul_109_11_n_472 & mul_109_11_n_441) | ((mul_109_11_n_441 & mul_109_11_n_560)
    | (mul_109_11_n_560 & mul_109_11_n_472)));
 assign mul_109_11_n_723 = (mul_109_11_n_441 ^ (mul_109_11_n_560 ^ mul_109_11_n_472));
 assign mul_109_11_n_720 = ((mul_109_11_n_458 & mul_109_11_n_620) | ((mul_109_11_n_620 & mul_109_11_n_447)
    | (mul_109_11_n_447 & mul_109_11_n_458)));
 assign mul_109_11_n_721 = (mul_109_11_n_620 ^ (mul_109_11_n_447 ^ mul_109_11_n_458));
 assign mul_109_11_n_718 = ((mul_109_11_n_463 & mul_109_11_n_593) | ((mul_109_11_n_593 & mul_109_11_n_426)
    | (mul_109_11_n_426 & mul_109_11_n_463)));
 assign mul_109_11_n_719 = (mul_109_11_n_593 ^ (mul_109_11_n_426 ^ mul_109_11_n_463));
 assign mul_109_11_n_716 = ((mul_109_11_n_536 & mul_109_11_n_629) | ((mul_109_11_n_629 & mul_109_11_n_422)
    | (mul_109_11_n_422 & mul_109_11_n_536)));
 assign mul_109_11_n_717 = (mul_109_11_n_629 ^ (mul_109_11_n_422 ^ mul_109_11_n_536));
 assign mul_109_11_n_715 = ~(mul_109_11_n_683 ^ mul_109_11_n_16);
 assign mul_109_11_n_714 = ~(mul_109_11_n_685 ^ mul_109_11_n_684);
 assign mul_109_11_n_712 = (mul_109_11_n_613 & mul_109_11_n_461);
 assign mul_109_11_n_713 = (mul_109_11_n_613 ^ mul_109_11_n_461);
 assign mul_109_11_n_710 = (mul_109_11_n_603 & mul_109_11_n_608);
 assign mul_109_11_n_711 = (mul_109_11_n_603 ^ mul_109_11_n_608);
 assign mul_109_11_n_708 = (mul_109_11_n_605 & mul_109_11_n_456);
 assign mul_109_11_n_709 = (mul_109_11_n_605 ^ mul_109_11_n_456);
 assign mul_109_11_n_706 = (mul_109_11_n_476 & mul_109_11_n_601);
 assign mul_109_11_n_707 = (mul_109_11_n_476 ^ mul_109_11_n_601);
 assign mul_109_11_n_704 = (mul_109_11_n_468 & mul_109_11_n_606);
 assign mul_109_11_n_705 = (mul_109_11_n_468 ^ mul_109_11_n_606);
 assign mul_109_11_n_702 = (mul_109_11_n_474 & mul_109_11_n_602);
 assign mul_109_11_n_703 = (mul_109_11_n_474 ^ mul_109_11_n_602);
 assign mul_109_11_n_700 = (mul_109_11_n_538 & mul_109_11_n_672);
 assign mul_109_11_n_701 = (mul_109_11_n_538 ^ mul_109_11_n_672);
 assign mul_109_11_n_698 = (mul_109_11_n_607 & mul_109_11_n_464);
 assign mul_109_11_n_699 = (mul_109_11_n_607 ^ mul_109_11_n_464);
 assign mul_109_11_n_696 = (mul_109_11_n_604 & mul_109_11_n_612);
 assign mul_109_11_n_697 = (mul_109_11_n_604 ^ mul_109_11_n_612);
 assign mul_109_11_n_694 = (mul_109_11_n_537 & mul_109_11_n_597);
 assign mul_109_11_n_695 = (mul_109_11_n_537 ^ mul_109_11_n_597);
 assign mul_109_11_n_692 = (mul_109_11_n_460 & mul_109_11_n_465);
 assign mul_109_11_n_693 = (mul_109_11_n_460 ^ mul_109_11_n_465);
 assign mul_109_11_n_690 = (mul_109_11_n_459 & mul_109_11_n_475);
 assign mul_109_11_n_691 = (mul_109_11_n_459 ^ mul_109_11_n_475);
 assign mul_109_11_n_688 = (mul_109_11_n_462 & mul_109_11_n_469);
 assign mul_109_11_n_689 = (mul_109_11_n_462 ^ mul_109_11_n_469);
 assign mul_109_11_n_686 = (mul_109_11_n_467 & mul_109_11_n_534);
 assign mul_109_11_n_687 = (mul_109_11_n_467 ^ mul_109_11_n_534);
 assign mul_109_11_n_685 = ~(mul_109_11_n_546 ^ mul_109_11_n_15);
 assign mul_109_11_n_684 = ~(mul_109_11_n_477 ^ mul_109_11_n_614);
 assign mul_109_11_n_683 = ~(mul_109_11_n_677 ^ mul_109_11_n_479);
 assign mul_109_11_n_682 = ~(mul_109_11_n_17 ^ mul_109_11_n_547);
 assign {out1[1]} = ~(mul_109_11_n_680 | (mul_109_11_n_548 & mul_109_11_n_329));
 assign mul_109_11_n_679 = ~((mul_109_11_n_412 & mul_109_11_n_276) | (mul_109_11_n_392 & mul_109_11_n_250));
 assign mul_109_11_n_678 = ~(mul_109_11_n_402 & (n_1448 & (mul_109_11_n_56 | mul_109_11_n_38)));
 assign mul_109_11_n_677 = ~((mul_109_11_n_14 | mul_109_11_n_303) & (mul_109_11_n_252 | mul_109_11_n_246));
 assign mul_109_11_n_676 = ~((mul_109_11_n_410 & mul_109_11_n_178) | (mul_109_11_n_391 & mul_109_11_n_81));
 assign mul_109_11_n_675 = ~((mul_109_11_n_408 & mul_109_11_n_107) | (mul_109_11_n_389 & mul_109_11_n_73));
 assign mul_109_11_n_674 = ~((mul_109_11_n_405 | mul_109_11_n_183) & (mul_109_11_n_257 | mul_109_11_n_212));
 assign mul_109_11_n_673 = ~((mul_109_11_n_13 | mul_109_11_n_301) & (mul_109_11_n_256 | mul_109_11_n_318));
 assign mul_109_11_n_670 = ~((mul_109_11_n_409 | mul_109_11_n_207) & (mul_109_11_n_263 | mul_109_11_n_192));
 assign mul_109_11_n_669 = ~((mul_109_11_n_409 | mul_109_11_n_192) & (mul_109_11_n_263 | mul_109_11_n_191));
 assign mul_109_11_n_668 = ~((mul_109_11_n_409 | mul_109_11_n_223) & (mul_109_11_n_263 | mul_109_11_n_207));
 assign mul_109_11_n_667 = ~((mul_109_11_n_406 | mul_109_11_n_105) & (mul_109_11_n_258 | mul_109_11_n_118));
 assign mul_109_11_n_663 = ~((mul_109_11_n_14 | mul_109_11_n_366) & (mul_109_11_n_252 | mul_109_11_n_303));
 assign mul_109_11_n_660 = ~((mul_109_11_n_407 | mul_109_11_n_94) & (mul_109_11_n_261 | mul_109_11_n_106));
 assign mul_109_11_n_659 = ~((mul_109_11_n_407 | mul_109_11_n_100) & (mul_109_11_n_261 | mul_109_11_n_92));
 assign mul_109_11_n_658 = ~((mul_109_11_n_407 | mul_109_11_n_75) & (mul_109_11_n_261 | mul_109_11_n_111));
 assign mul_109_11_n_657 = ~((mul_109_11_n_407 | mul_109_11_n_92) & (mul_109_11_n_261 | mul_109_11_n_93));
 assign mul_109_11_n_656 = ~((mul_109_11_n_407 | mul_109_11_n_101) & (mul_109_11_n_261 | mul_109_11_n_100));
 assign mul_109_11_n_655 = ~((mul_109_11_n_407 | mul_109_11_n_111) & (mul_109_11_n_261 | mul_109_11_n_101));
 assign mul_109_11_n_654 = ~((mul_109_11_n_407 | mul_109_11_n_93) & (mul_109_11_n_261 | mul_109_11_n_95));
 assign mul_109_11_n_653 = ~((mul_109_11_n_407 | mul_109_11_n_95) & (mul_109_11_n_261 | mul_109_11_n_94));
 assign mul_109_11_n_652 = ~((mul_109_11_n_406 | mul_109_11_n_164) & (mul_109_11_n_258 | mul_109_11_n_165));
 assign mul_109_11_n_651 = ~((mul_109_11_n_406 | mul_109_11_n_196) & (mul_109_11_n_258 | mul_109_11_n_87));
 assign mul_109_11_n_650 = ~((mul_109_11_n_406 | mul_109_11_n_86) & (mul_109_11_n_258 | mul_109_11_n_372));
 assign mul_109_11_n_649 = ~((mul_109_11_n_406 | mul_109_11_n_118) & (mul_109_11_n_258 | mul_109_11_n_117));
 assign mul_109_11_n_680 = ~(mul_109_11_n_548 | mul_109_11_n_329);
 assign mul_109_11_n_648 = ~((mul_109_11_n_406 | mul_109_11_n_77) & (mul_109_11_n_258 | mul_109_11_n_105));
 assign mul_109_11_n_647 = ~((mul_109_11_n_406 | mul_109_11_n_143) & (mul_109_11_n_258 | mul_109_11_n_164));
 assign mul_109_11_n_646 = ~((mul_109_11_n_406 | mul_109_11_n_195) & (mul_109_11_n_258 | mul_109_11_n_196));
 assign mul_109_11_n_645 = ~((mul_109_11_n_406 | mul_109_11_n_87) & (mul_109_11_n_258 | mul_109_11_n_86));
 assign mul_109_11_n_644 = ~((mul_109_11_n_406 | mul_109_11_n_142) & (mul_109_11_n_258 | mul_109_11_n_143));
 assign mul_109_11_n_643 = ~((mul_109_11_n_406 | mul_109_11_n_165) & (mul_109_11_n_258 | mul_109_11_n_195));
 assign mul_109_11_n_642 = ~((mul_109_11_n_406 | mul_109_11_n_129) & (mul_109_11_n_258 | mul_109_11_n_128));
 assign mul_109_11_n_641 = ~((mul_109_11_n_406 | mul_109_11_n_128) & (mul_109_11_n_258 | mul_109_11_n_142));
 assign mul_109_11_n_640 = ~((mul_109_11_n_406 | mul_109_11_n_117) & (mul_109_11_n_258 | mul_109_11_n_129));
 assign mul_109_11_n_639 = ~((mul_109_11_n_411 | mul_109_11_n_282) & (mul_109_11_n_264 | mul_109_11_n_275));
 assign mul_109_11_n_638 = ~((mul_109_11_n_405 | mul_109_11_n_139) & (mul_109_11_n_257 | mul_109_11_n_158));
 assign mul_109_11_n_637 = ~((mul_109_11_n_405 | mul_109_11_n_138) & (mul_109_11_n_257 | mul_109_11_n_139));
 assign mul_109_11_n_636 = ~((mul_109_11_n_405 | mul_109_11_n_151) & (mul_109_11_n_257 | mul_109_11_n_149));
 assign mul_109_11_n_635 = ~((mul_109_11_n_405 | mul_109_11_n_127) & (mul_109_11_n_257 | mul_109_11_n_138));
 assign mul_109_11_n_634 = ~((mul_109_11_n_405 | mul_109_11_n_157) & (mul_109_11_n_257 | mul_109_11_n_184));
 assign mul_109_11_n_633 = ~((mul_109_11_n_405 | mul_109_11_n_272) & (mul_109_11_n_257 | mul_109_11_n_296));
 assign mul_109_11_n_632 = ~((mul_109_11_n_405 | mul_109_11_n_184) & (mul_109_11_n_257 | mul_109_11_n_183));
 assign mul_109_11_n_631 = ~((mul_109_11_n_405 | mul_109_11_n_149) & (mul_109_11_n_257 | mul_109_11_n_271));
 assign mul_109_11_n_629 = ~((mul_109_11_n_405 | mul_109_11_n_213) & (mul_109_11_n_257 | mul_109_11_n_151));
 assign mul_109_11_n_628 = ~((mul_109_11_n_405 | mul_109_11_n_126) & (mul_109_11_n_257 | mul_109_11_n_127));
 assign mul_109_11_n_627 = ~((mul_109_11_n_405 | mul_109_11_n_119) & (mul_109_11_n_257 | mul_109_11_n_126));
 assign mul_109_11_n_626 = ~((mul_109_11_n_405 | mul_109_11_n_76) & (mul_109_11_n_257 | mul_109_11_n_119));
 assign mul_109_11_n_625 = ~((mul_109_11_n_405 | mul_109_11_n_271) & (mul_109_11_n_257 | mul_109_11_n_272));
 assign mul_109_11_n_624 = ~((mul_109_11_n_405 | mul_109_11_n_212) & (mul_109_11_n_257 | mul_109_11_n_213));
 assign mul_109_11_n_623 = ~((mul_109_11_n_405 | mul_109_11_n_158) & (mul_109_11_n_257 | mul_109_11_n_157));
 assign mul_109_11_n_622 = ~((mul_109_11_n_411 | mul_109_11_n_227) & (mul_109_11_n_264 | mul_109_11_n_282));
 assign mul_109_11_n_621 = ~((mul_109_11_n_13 | mul_109_11_n_278) & (mul_109_11_n_256 | mul_109_11_n_279));
 assign mul_109_11_n_620 = ~((mul_109_11_n_13 | mul_109_11_n_279) & (mul_109_11_n_256 | mul_109_11_n_302));
 assign mul_109_11_n_619 = ~((mul_109_11_n_409 | mul_109_11_n_191) & (mul_109_11_n_263 | mul_109_11_n_177));
 assign mul_109_11_n_618 = ~((mul_109_11_n_13 | mul_109_11_n_154) & (mul_109_11_n_256 | mul_109_11_n_171));
 assign mul_109_11_n_617 = ~((mul_109_11_n_13 | mul_109_11_n_153) & (mul_109_11_n_256 | mul_109_11_n_154));
 assign mul_109_11_n_616 = ~((mul_109_11_n_13 | mul_109_11_n_85) & (mul_109_11_n_256 | mul_109_11_n_334));
 assign mul_109_11_n_614 = ((mul_109_11_n_256 | mul_109_11_n_226) & (mul_109_11_n_13 | mul_109_11_n_318));
 assign mul_109_11_n_615 = ~((mul_109_11_n_14 | mul_109_11_n_69) & (mul_109_11_n_252 | mul_109_11_n_159));
 assign mul_109_11_n_606 = ~((mul_109_11_n_13 | mul_109_11_n_302) & (mul_109_11_n_256 | mul_109_11_n_301));
 assign mul_109_11_n_604 = ~((mul_109_11_n_14 | mul_109_11_n_277) & (mul_109_11_n_252 | mul_109_11_n_375));
 assign mul_109_11_n_603 = ~((mul_109_11_n_14 | mul_109_11_n_134) & (mul_109_11_n_252 | mul_109_11_n_120));
 assign mul_109_11_n_602 = ~((mul_109_11_n_14 | mul_109_11_n_214) & (mul_109_11_n_252 | mul_109_11_n_215));
 assign mul_109_11_n_601 = ~((mul_109_11_n_14 | mul_109_11_n_193) & (mul_109_11_n_252 | mul_109_11_n_194));
 assign mul_109_11_n_600 = ~((mul_109_11_n_13 | mul_109_11_n_334) & (mul_109_11_n_256 | mul_109_11_n_322));
 assign mul_109_11_n_599 = ~((mul_109_11_n_14 | mul_109_11_n_297) & (mul_109_11_n_252 | mul_109_11_n_313));
 assign mul_109_11_n_598 = ~((mul_109_11_n_14 | mul_109_11_n_280) & (mul_109_11_n_252 | mul_109_11_n_298));
 assign mul_109_11_n_596 = ~((mul_109_11_n_13 | mul_109_11_n_84) & (mul_109_11_n_256 | mul_109_11_n_123));
 assign mul_109_11_n_594 = ~((mul_109_11_n_13 | mul_109_11_n_200) & (mul_109_11_n_256 | mul_109_11_n_221));
 assign mul_109_11_n_592 = ~((mul_109_11_n_13 | mul_109_11_n_322) & (mul_109_11_n_256 | mul_109_11_n_278));
 assign mul_109_11_n_582 = ~((mul_109_11_n_13 | mul_109_11_n_171) & (mul_109_11_n_256 | mul_109_11_n_172));
 assign mul_109_11_n_580 = ~((mul_109_11_n_13 | mul_109_11_n_136) & (mul_109_11_n_256 | mul_109_11_n_153));
 assign mul_109_11_n_579 = ~((mul_109_11_n_13 | mul_109_11_n_199) & (mul_109_11_n_256 | mul_109_11_n_200));
 assign mul_109_11_n_578 = ~((mul_109_11_n_14 | mul_109_11_n_298) & (mul_109_11_n_252 | mul_109_11_n_297));
 assign mul_109_11_n_577 = ~((mul_109_11_n_14 | mul_109_11_n_353) & (mul_109_11_n_252 | mul_109_11_n_352));
 assign mul_109_11_n_576 = ~((mul_109_11_n_14 | mul_109_11_n_281) & (mul_109_11_n_252 | mul_109_11_n_280));
 assign mul_109_11_n_575 = ~((mul_109_11_n_13 | mul_109_11_n_221) & (mul_109_11_n_256 | mul_109_11_n_85));
 assign mul_109_11_n_574 = ~((mul_109_11_n_14 | mul_109_11_n_375) & (mul_109_11_n_252 | mul_109_11_n_281));
 assign mul_109_11_n_573 = ~((mul_109_11_n_14 | mul_109_11_n_352) & (mul_109_11_n_252 | mul_109_11_n_367));
 assign mul_109_11_n_572 = ~((mul_109_11_n_14 | mul_109_11_n_328) & (mul_109_11_n_252 | mul_109_11_n_340));
 assign mul_109_11_n_571 = ~((mul_109_11_n_14 | mul_109_11_n_340) & (mul_109_11_n_252 | mul_109_11_n_341));
 assign mul_109_11_n_570 = ~((mul_109_11_n_14 | mul_109_11_n_120) & (mul_109_11_n_252 | mul_109_11_n_277));
 assign mul_109_11_n_569 = ~((mul_109_11_n_14 | mul_109_11_n_327) & (mul_109_11_n_252 | mul_109_11_n_328));
 assign mul_109_11_n_567 = ~((mul_109_11_n_14 | mul_109_11_n_312) & (mul_109_11_n_252 | mul_109_11_n_327));
 assign mul_109_11_n_566 = ~((mul_109_11_n_14 | mul_109_11_n_215) & (mul_109_11_n_252 | mul_109_11_n_134));
 assign mul_109_11_n_565 = ~((mul_109_11_n_13 | mul_109_11_n_137) & (mul_109_11_n_256 | mul_109_11_n_136));
 assign mul_109_11_n_564 = ~((mul_109_11_n_14 | mul_109_11_n_194) & (mul_109_11_n_252 | mul_109_11_n_214));
 assign mul_109_11_n_563 = ~((mul_109_11_n_14 | mul_109_11_n_341) & (mul_109_11_n_252 | mul_109_11_n_353));
 assign mul_109_11_n_561 = ~((mul_109_11_n_14 | mul_109_11_n_174) & (mul_109_11_n_252 | mul_109_11_n_173));
 assign mul_109_11_n_560 = ~((mul_109_11_n_14 | mul_109_11_n_313) & (mul_109_11_n_252 | mul_109_11_n_312));
 assign mul_109_11_n_559 = ~((mul_109_11_n_14 | mul_109_11_n_173) & (mul_109_11_n_252 | mul_109_11_n_193));
 assign mul_109_11_n_558 = ~((mul_109_11_n_14 | mul_109_11_n_367) & (mul_109_11_n_252 | mul_109_11_n_366));
 assign mul_109_11_n_556 = ~((mul_109_11_n_14 | mul_109_11_n_159) & (mul_109_11_n_252 | mul_109_11_n_174));
 assign mul_109_11_n_555 = ~((mul_109_11_n_13 | mul_109_11_n_123) & (mul_109_11_n_256 | mul_109_11_n_137));
 assign mul_109_11_n_549 = ~((mul_109_11_n_13 | mul_109_11_n_172) & (mul_109_11_n_256 | mul_109_11_n_199));
 assign mul_109_11_n_545 = ~((mul_109_11_n_266 | (mul_109_11_n_225 | mul_109_11_n_0)) & (mul_109_11_n_265
    | mul_109_11_n_232));
 assign mul_109_11_n_544 = ~((mul_109_11_n_384 | mul_109_11_n_170) & (mul_109_11_n_190 | mul_109_11_n_26));
 assign mul_109_11_n_543 = ~((mul_109_11_n_387 | mul_109_11_n_109) & (mul_109_11_n_262 | mul_109_11_n_74));
 assign mul_109_11_n_542 = ~((mul_109_11_n_386 | mul_109_11_n_148) & (mul_109_11_n_260 | mul_109_11_n_78));
 assign mul_109_11_n_541 = ~((mul_109_11_n_385 | mul_109_11_n_206) & (mul_109_11_n_259 | mul_109_11_n_83));
 assign mul_109_11_n_540 = ~((mul_109_11_n_384 | mul_109_11_n_374) & (mul_109_11_n_347 | mul_109_11_n_26));
 assign mul_109_11_n_539 = ~((mul_109_11_n_384 | mul_109_11_n_365) & (mul_109_11_n_295 | mul_109_11_n_26));
 assign mul_109_11_n_538 = ~((mul_109_11_n_384 | mul_109_11_n_208) & (mul_109_11_n_209 | mul_109_11_n_26));
 assign mul_109_11_n_537 = ~((mul_109_11_n_384 | mul_109_11_n_190) & (mul_109_11_n_189 | mul_109_11_n_26));
 assign mul_109_11_n_536 = ~((mul_109_11_n_384 | mul_109_11_n_370) & (mul_109_11_n_294 | mul_109_11_n_26));
 assign mul_109_11_n_535 = ~((mul_109_11_n_385 | mul_109_11_n_104) & (mul_109_11_n_259 | mul_109_11_n_103));
 assign mul_109_11_n_534 = ~((mul_109_11_n_384 | mul_109_11_n_108) & (mul_109_11_n_102 | mul_109_11_n_26));
 assign mul_109_11_n_533 = ~((mul_109_11_n_384 | mul_109_11_n_361) & (mul_109_11_n_161 | mul_109_11_n_26));
 assign mul_109_11_n_532 = ~((mul_109_11_n_384 | mul_109_11_n_161) & (mul_109_11_n_267 | mul_109_11_n_26));
 assign mul_109_11_n_531 = ~((mul_109_11_n_384 | mul_109_11_n_294) & (mul_109_11_n_365 | mul_109_11_n_26));
 assign mul_109_11_n_530 = ~((mul_109_11_n_384 | mul_109_11_n_209) & (mul_109_11_n_108 | mul_109_11_n_26));
 assign mul_109_11_n_529 = ~((mul_109_11_n_384 | mul_109_11_n_333) & (mul_109_11_n_332 | mul_109_11_n_26));
 assign mul_109_11_n_528 = ~((mul_109_11_n_384 | mul_109_11_n_332) & (mul_109_11_n_345 | mul_109_11_n_26));
 assign mul_109_11_n_527 = ~((mul_109_11_n_384 | mul_109_11_n_344) & (mul_109_11_n_356 | mul_109_11_n_26));
 assign mul_109_11_n_526 = ~((mul_109_11_n_384 | mul_109_11_n_317) & (mul_109_11_n_333 | mul_109_11_n_26));
 assign mul_109_11_n_525 = ~((mul_109_11_n_384 | mul_109_11_n_345) & (mul_109_11_n_344 | mul_109_11_n_26));
 assign mul_109_11_n_524 = ~((mul_109_11_n_384 | mul_109_11_n_316) & (mul_109_11_n_317 | mul_109_11_n_26));
 assign mul_109_11_n_523 = ~((mul_109_11_n_384 | mul_109_11_n_189) & (mul_109_11_n_208 | mul_109_11_n_26));
 assign mul_109_11_n_522 = ~((mul_109_11_n_384 | mul_109_11_n_357) & (mul_109_11_n_371 | mul_109_11_n_26));
 assign mul_109_11_n_518 = ~((mul_109_11_n_384 | mul_109_11_n_102) & (mul_109_11_n_361 | mul_109_11_n_26));
 assign mul_109_11_n_517 = ~((mul_109_11_n_384 | mul_109_11_n_304) & (mul_109_11_n_316 | mul_109_11_n_26));
 assign mul_109_11_n_516 = ~((mul_109_11_n_384 | mul_109_11_n_371) & (mul_109_11_n_370 | mul_109_11_n_26));
 assign mul_109_11_n_515 = ~((mul_109_11_n_384 | mul_109_11_n_295) & (mul_109_11_n_374 | mul_109_11_n_26));
 assign mul_109_11_n_514 = ~((mul_109_11_n_384 | mul_109_11_n_305) & (mul_109_11_n_304 | mul_109_11_n_26));
 assign mul_109_11_n_513 = ~((mul_109_11_n_384 | mul_109_11_n_287) & (mul_109_11_n_305 | mul_109_11_n_26));
 assign mul_109_11_n_512 = ~((mul_109_11_n_384 | mul_109_11_n_356) & (mul_109_11_n_357 | mul_109_11_n_26));
 assign mul_109_11_n_511 = ~((mul_109_11_n_387 | mul_109_11_n_121) & (mul_109_11_n_262 | mul_109_11_n_109));
 assign mul_109_11_n_510 = ~((mul_109_11_n_387 | mul_109_11_n_122) & (mul_109_11_n_262 | mul_109_11_n_121));
 assign mul_109_11_n_509 = ~((mul_109_11_n_387 | mul_109_11_n_140) & (mul_109_11_n_262 | mul_109_11_n_132));
 assign mul_109_11_n_508 = ~((mul_109_11_n_387 | mul_109_11_n_132) & (mul_109_11_n_262 | mul_109_11_n_133));
 assign mul_109_11_n_507 = ~((mul_109_11_n_387 | mul_109_11_n_237) & (mul_109_11_n_262 | mul_109_11_n_140));
 assign mul_109_11_n_506 = ~((mul_109_11_n_387 | mul_109_11_n_133) & (mul_109_11_n_262 | mul_109_11_n_122));
 assign mul_109_11_n_505 = ~((mul_109_11_n_386 | mul_109_11_n_82) & (mul_109_11_n_260 | mul_109_11_n_88));
 assign mul_109_11_n_504 = ~((mul_109_11_n_386 | mul_109_11_n_88) & (mul_109_11_n_260 | mul_109_11_n_89));
 assign mul_109_11_n_503 = ~((mul_109_11_n_386 | mul_109_11_n_124) & (mul_109_11_n_260 | mul_109_11_n_148));
 assign mul_109_11_n_502 = ~((mul_109_11_n_386 | mul_109_11_n_99) & (mul_109_11_n_260 | mul_109_11_n_98));
 assign mul_109_11_n_501 = ~((mul_109_11_n_386 | mul_109_11_n_98) & (mul_109_11_n_260 | mul_109_11_n_113));
 assign mul_109_11_n_500 = ~((mul_109_11_n_386 | mul_109_11_n_90) & (mul_109_11_n_260 | mul_109_11_n_99));
 assign mul_109_11_n_499 = ~((mul_109_11_n_386 | mul_109_11_n_89) & (mul_109_11_n_260 | mul_109_11_n_90));
 assign mul_109_11_n_498 = ~((mul_109_11_n_386 | mul_109_11_n_113) & (mul_109_11_n_260 | mul_109_11_n_114));
 assign mul_109_11_n_497 = ~((mul_109_11_n_386 | mul_109_11_n_125) & (mul_109_11_n_260 | mul_109_11_n_124));
 assign mul_109_11_n_496 = ~((mul_109_11_n_384 | mul_109_11_n_288) & (mul_109_11_n_287 | mul_109_11_n_26));
 assign mul_109_11_n_495 = ~((mul_109_11_n_386 | mul_109_11_n_114) & (mul_109_11_n_260 | mul_109_11_n_125));
 assign mul_109_11_n_494 = ~((mul_109_11_n_385 | mul_109_11_n_79) & (mul_109_11_n_259 | mul_109_11_n_96));
 assign mul_109_11_n_493 = ~((mul_109_11_n_384 | mul_109_11_n_267) & (mul_109_11_n_268 | mul_109_11_n_26));
 assign mul_109_11_n_492 = ~((mul_109_11_n_385 | mul_109_11_n_131) & (mul_109_11_n_259 | mul_109_11_n_130));
 assign mul_109_11_n_491 = ~((mul_109_11_n_385 | mul_109_11_n_168) & (mul_109_11_n_259 | mul_109_11_n_206));
 assign mul_109_11_n_490 = ~((mul_109_11_n_385 | mul_109_11_n_144) & (mul_109_11_n_259 | mul_109_11_n_167));
 assign mul_109_11_n_489 = ~((mul_109_11_n_385 | mul_109_11_n_115) & (mul_109_11_n_259 | mul_109_11_n_131));
 assign mul_109_11_n_488 = ~((mul_109_11_n_385 | mul_109_11_n_145) & (mul_109_11_n_259 | mul_109_11_n_144));
 assign mul_109_11_n_487 = ~((mul_109_11_n_385 | mul_109_11_n_130) & (mul_109_11_n_259 | mul_109_11_n_145));
 assign mul_109_11_n_486 = ~((mul_109_11_n_385 | mul_109_11_n_116) & (mul_109_11_n_259 | mul_109_11_n_115));
 assign mul_109_11_n_485 = ~((mul_109_11_n_385 | mul_109_11_n_96) & (mul_109_11_n_259 | mul_109_11_n_104));
 assign mul_109_11_n_484 = ~((mul_109_11_n_385 | mul_109_11_n_103) & (mul_109_11_n_259 | mul_109_11_n_116));
 assign mul_109_11_n_483 = ~((mul_109_11_n_385 | mul_109_11_n_167) & (mul_109_11_n_259 | mul_109_11_n_168));
 assign mul_109_11_n_482 = ~((mul_109_11_n_384 | mul_109_11_n_268) & (mul_109_11_n_288 | mul_109_11_n_26));
 assign mul_109_11_n_481 = ~((mul_109_11_n_12 | mul_109_11_n_210) & (mul_109_11_n_255 | mul_109_11_n_211));
 assign mul_109_11_n_479 = ~((mul_109_11_n_12 | mul_109_11_n_335) & (mul_109_11_n_255 | mul_109_11_n_228));
 assign mul_109_11_n_475 = ~((mul_109_11_n_12 | mul_109_11_n_306) & (mul_109_11_n_255 | mul_109_11_n_307));
 assign mul_109_11_n_469 = ~((mul_109_11_n_12 | mul_109_11_n_360) & (mul_109_11_n_255 | mul_109_11_n_346));
 assign mul_109_11_n_468 = ~((mul_109_11_n_12 | mul_109_11_n_321) & (mul_109_11_n_255 | mul_109_11_n_320));
 assign mul_109_11_n_465 = ~((mul_109_11_n_12 | mul_109_11_n_286) & (mul_109_11_n_255 | mul_109_11_n_285));
 assign mul_109_11_n_449 = ~((mul_109_11_n_12 | mul_109_11_n_346) & (mul_109_11_n_255 | mul_109_11_n_286));
 assign mul_109_11_n_448 = ~((mul_109_11_n_12 | mul_109_11_n_285) & (mul_109_11_n_255 | mul_109_11_n_306));
 assign mul_109_11_n_447 = ~((mul_109_11_n_12 | mul_109_11_n_307) & (mul_109_11_n_255 | mul_109_11_n_321));
 assign mul_109_11_n_446 = ~((mul_109_11_n_12 | mul_109_11_n_211) & (mul_109_11_n_255 | mul_109_11_n_110));
 assign mul_109_11_n_444 = ~((mul_109_11_n_12 | mul_109_11_n_72) & (mul_109_11_n_255 | mul_109_11_n_135));
 assign mul_109_11_n_441 = ~((mul_109_11_n_12 | mul_109_11_n_110) & (mul_109_11_n_255 | mul_109_11_n_112));
 assign mul_109_11_n_437 = ~((mul_109_11_n_12 | mul_109_11_n_135) & (mul_109_11_n_255 | mul_109_11_n_147));
 assign mul_109_11_n_436 = ~((mul_109_11_n_12 | mul_109_11_n_147) & (mul_109_11_n_255 | mul_109_11_n_146));
 assign mul_109_11_n_431 = ~((mul_109_11_n_12 | mul_109_11_n_146) & (mul_109_11_n_255 | mul_109_11_n_162));
 assign mul_109_11_n_426 = ~((mul_109_11_n_12 | mul_109_11_n_112) & (mul_109_11_n_255 | mul_109_11_n_360));
 assign mul_109_11_n_425 = ~((mul_109_11_n_12 | mul_109_11_n_162) & (mul_109_11_n_255 | mul_109_11_n_163));
 assign mul_109_11_n_423 = ~((mul_109_11_n_12 | mul_109_11_n_187) & (mul_109_11_n_255 | mul_109_11_n_210));
 assign mul_109_11_n_420 = ~((mul_109_11_n_12 | mul_109_11_n_163) & (mul_109_11_n_255 | mul_109_11_n_188));
 assign mul_109_11_n_416 = ~((mul_109_11_n_12 | mul_109_11_n_188) & (mul_109_11_n_255 | mul_109_11_n_187));
 assign mul_109_11_n_413 = ~((mul_109_11_n_12 | mul_109_11_n_320) & (mul_109_11_n_255 | mul_109_11_n_335));
 assign mul_109_11_n_412 = ~mul_109_11_n_411;
 assign mul_109_11_n_410 = ~mul_109_11_n_409;
 assign mul_109_11_n_408 = ~mul_109_11_n_407;
 assign mul_109_11_n_411 = ~(mul_109_11_n_264 & mul_109_11_n_230);
 assign mul_109_11_n_409 = ~(mul_109_11_n_263 & mul_109_11_n_231);
 assign mul_109_11_n_407 = ~(mul_109_11_n_261 & mul_109_11_n_236);
 assign mul_109_11_n_406 = (mul_109_11_n_388 | mul_109_11_n_240);
 assign mul_109_11_n_405 = (mul_109_11_n_390 | mul_109_11_n_241);
 assign mul_109_11_n_404 = (mul_109_11_n_393 | mul_109_11_n_245);
 assign mul_109_11_n_401 = ~(mul_109_11_n_258 | mul_109_11_n_38);
 assign mul_109_11_n_400 = ~(mul_109_11_n_256 | mul_109_11_n_38);
 assign mul_109_11_n_399 = ~(mul_109_11_n_252 | mul_109_11_n_38);
 assign mul_109_11_n_398 = ~(mul_109_11_n_257 | mul_109_11_n_38);
 assign mul_109_11_n_397 = ~(mul_109_11_n_261 | mul_109_11_n_38);
 assign mul_109_11_n_396 = ~(mul_109_11_n_263 | mul_109_11_n_38);
 assign mul_109_11_n_394 = ~(mul_109_11_n_264 | mul_109_11_n_38);
 assign mul_109_11_n_392 = ~mul_109_11_n_264;
 assign mul_109_11_n_391 = ~mul_109_11_n_263;
 assign mul_109_11_n_390 = ~mul_109_11_n_257;
 assign mul_109_11_n_389 = ~mul_109_11_n_261;
 assign mul_109_11_n_388 = ~mul_109_11_n_258;
 assign mul_109_11_n_383 = ~mul_109_11_n_384;
 assign mul_109_11_n_382 = ~(mul_109_11_n_265 | mul_109_11_n_38);
 assign mul_109_11_n_387 = ~(mul_109_11_n_262 & mul_109_11_n_235);
 assign mul_109_11_n_386 = ~(mul_109_11_n_260 & mul_109_11_n_238);
 assign mul_109_11_n_385 = ~(mul_109_11_n_259 & mul_109_11_n_239);
 assign mul_109_11_n_380 = ~(mul_109_11_n_260 | mul_109_11_n_38);
 assign mul_109_11_n_379 = ~(mul_109_11_n_259 | mul_109_11_n_38);
 assign mul_109_11_n_378 = ~(mul_109_11_n_255 | mul_109_11_n_38);
 assign mul_109_11_n_377 = ~(mul_109_11_n_262 | mul_109_11_n_38);
 assign mul_109_11_n_348 = ~mul_109_11_n_347;
 assign mul_109_11_n_276 = ~mul_109_11_n_275;
 assign mul_109_11_n_266 = ~mul_109_11_n_265;
 assign mul_109_11_n_236 = ~((mul_109_11_n_28 & ~n_1457) | (n_1456 & n_1457));
 assign mul_109_11_n_235 = ~((mul_109_11_n_31 & ~n_1455) | (n_1454 & n_1455));
 assign mul_109_11_n_231 = ~((mul_109_11_n_52 & ~n_1453) | (n_1452 & n_1453));
 assign mul_109_11_n_230 = ~((mul_109_11_n_56 & ~n_1451) | (n_1450 & n_1451));
 assign mul_109_11_n_225 = ~(n_1448 ^ n_1449);
 assign mul_109_11_n_265 = ~(n_1449 ^ n_1450);
 assign mul_109_11_n_264 = ((mul_109_11_n_52 & ~n_1451) | (n_1452 & n_1451));
 assign mul_109_11_n_263 = ~(n_1453 ^ n_1454);
 assign mul_109_11_n_262 = ~(n_1455 ^ n_1456);
 assign mul_109_11_n_261 = ~(n_1457 ^ n_1458);
 assign mul_109_11_n_178 = ~mul_109_11_n_177;
 assign mul_109_11_n_170 = ~mul_109_11_n_169;
 assign mul_109_11_n_107 = ~mul_109_11_n_106;
 assign mul_109_11_n_65 = ~(mul_109_11_n_19 & mul_109_11_n_38);
 assign mul_109_11_n_64 = ~(mul_109_11_n_28 & mul_109_11_n_38);
 assign mul_109_11_n_63 = ~(mul_109_11_n_41 & mul_109_11_n_38);
 assign mul_109_11_n_62 = ~(mul_109_11_n_25 & mul_109_11_n_38);
 assign mul_109_11_n_61 = ~(mul_109_11_n_39 & mul_109_11_n_38);
 assign {out1[0]} = ~(mul_109_11_n_26 | mul_109_11_n_38);
 assign mul_109_11_n_56 = ~n_1450;
 assign mul_109_11_n_52 = ~n_1452;
 assign mul_109_11_n_43 = ~n_1458;
 assign mul_109_11_n_31 = ~n_1454;
 assign mul_109_11_n_28 = ~n_1456;
 assign mul_109_11_n_17 = ~(~(mul_109_11_n_406 | mul_109_11_n_372) | (mul_109_11_n_388 & mul_109_11_n_234));
 assign mul_109_11_n_16 = ~(~(mul_109_11_n_405 | mul_109_11_n_296) | (mul_109_11_n_390 & mul_109_11_n_224));
 assign mul_109_11_n_15 = ~(~(mul_109_11_n_404 | mul_109_11_n_364) | (mul_109_11_n_393 & mul_109_11_n_233));
 assign mul_109_11_n_14 = ~(mul_109_11_n_252 & ~mul_109_11_n_247);
 assign mul_109_11_n_13 = ~(mul_109_11_n_256 & ~mul_109_11_n_242);
 assign mul_109_11_n_12 = ~(mul_109_11_n_255 & ~n_1493);
 assign mul_109_11_n_3 = ~(mul_109_11_n_52 & ~n_1451);
 assign mul_109_11_n_2 = ~(mul_109_11_n_43 & ~n_1457);
 assign mul_109_11_n_1 = ~(mul_109_11_n_31 & ~n_1453);
 assign n_1479 = ~(csa_tree_add_64_2_groupi_n_8 ^ csa_tree_add_64_2_groupi_n_64);
 assign n_1480 = ({in5[1]} ^ {in6[1]});
 assign n_1482 = ((n_1481 & ~csa_tree_add_71_2_groupi_n_54) | (csa_tree_add_71_2_groupi_n_119 & csa_tree_add_71_2_groupi_n_54));
 assign n_1481 = ~(csa_tree_add_71_2_groupi_n_116 | ~csa_tree_add_71_2_groupi_n_62);
 assign n_1483 = (csa_tree_add_71_2_groupi_n_57 ^ csa_tree_add_71_2_groupi_n_52);
 assign n_1484 = ~(csa_tree_add_71_2_groupi_n_109 ^ csa_tree_add_71_2_groupi_n_87);
 assign n_1486 = (csa_tree_add_71_2_groupi_n_103 ^ n_1485);
 assign n_1485 = ~(csa_tree_add_71_2_groupi_n_72 & csa_tree_add_71_2_groupi_n_64);
 assign n_1487 = (n_1488 ^ {in1[0]});
 assign n_1488 = ({in3[0]} ^ {in2[0]});
 assign n_1489 = ~(csa_tree_mul_77_11_groupi_n_14 & (n_1321 & ~n_1322));
 assign n_1490 = ((n_1500 & ~csa_tree_mul_77_11_groupi_n_12) | (csa_tree_mul_77_11_groupi_n_21 & csa_tree_mul_77_11_groupi_n_12));
 assign n_1491 = ((n_1306 & ~csa_tree_mul_77_11_groupi_n_13) | (csa_tree_mul_77_11_groupi_n_16 & csa_tree_mul_77_11_groupi_n_13));
 assign n_1492 = ~(csa_tree_add_106_2_groupi_n_45 & (n_1437 & ~n_1438));
 assign n_1493 = ~((n_81 & ~n_84) | (n_1185 & n_84));
 assign n_1494 = ~((n_1324 & ~n_104) | (n_1336 & n_104));
 assign n_1495 = ~(csa_tree_mul_77_11_groupi_n_549 ^ csa_tree_mul_77_11_groupi_n_6);
 assign n_1496 = ~(csa_tree_mul_77_11_groupi_n_451 ^ csa_tree_mul_77_11_groupi_n_492);
 assign n_1497 = ~(csa_tree_mul_77_11_groupi_n_409 ^ csa_tree_mul_77_11_groupi_n_416);
 assign n_1498 = (csa_tree_mul_77_11_groupi_n_570 ^ csa_tree_mul_77_11_groupi_n_9);
 assign n_1499 = ~(csa_tree_add_106_2_groupi_n_46 & (n_1446 & ~n_1447));
 assign n_1500 = ~(mul_74_11_n_501 ^ mul_74_11_n_498);
 assign n_1501 = ~(mul_74_11_n_482 ^ mul_74_11_n_459);
 assign n_1502 = ~(mul_74_11_n_452 ^ mul_74_11_n_472);
 assign n_1503 = ~(mul_74_11_n_442 ^ mul_74_11_n_437);
 assign n_1504 = (mul_74_11_n_326 ^ mul_74_11_n_218);
 assign n_1505 = (mul_74_11_n_284 ^ mul_74_11_n_241);
 assign n_1506 = ~(n_1292 & mul_74_11_n_47);
 assign n_1508 = (mul_74_11_n_169 & n_1507);
 assign n_1507 = ~((n_1482 & ~mul_74_11_n_44) | (mul_74_11_n_37 & mul_74_11_n_44));
 assign n_1510 = ~(n_1518 | n_1509);
 assign n_1509 = ~((n_1484 & ~n_1486) | (mul_74_11_n_30 & n_1486));
 assign n_1511 = ((n_1482 & ~n_1277) | (mul_74_11_n_37 & n_1277));
 assign n_1512 = ((n_1482 & ~n_1280) | (mul_74_11_n_37 & n_1280));
 assign n_1513 = ((n_1275 & ~mul_74_11_n_35) | (mul_74_11_n_39 & mul_74_11_n_35));
 assign n_1514 = ((n_1280 & ~mul_74_11_n_35) | (mul_74_11_n_40 & mul_74_11_n_35));
 assign n_1515 = ((n_1276 & ~mul_74_11_n_35) | (mul_74_11_n_50 & mul_74_11_n_35));
 assign n_1516 = ((n_1274 & ~mul_74_11_n_35) | (mul_74_11_n_51 & mul_74_11_n_35));
 assign n_1517 = ((n_1276 & ~mul_74_11_n_37) | (mul_74_11_n_50 & mul_74_11_n_37));
 assign n_1518 = (n_1292 ^ n_1486);
 assign n_1519 = ((n_1292 & ~mul_74_11_n_46) | (mul_74_11_n_35 & mul_74_11_n_46));
 assign n_1520 = ((n_1482 & ~n_1283) | (mul_74_11_n_37 & n_1283));
 assign n_1521 = ((n_1286 & ~mul_74_11_n_46) | (mul_74_11_n_45 & mul_74_11_n_46));
 assign n_1522 = ((mul_74_11_n_31 & ~n_1282) | (mul_74_11_n_30 & n_1282));
 assign n_1523 = ((n_1286 & ~n_1282) | (mul_74_11_n_45 & n_1282));
 assign n_1524 = ((n_1275 & ~mul_74_11_n_30) | (mul_74_11_n_39 & mul_74_11_n_30));
 assign n_1525 = ((n_1276 & ~mul_74_11_n_30) | (mul_74_11_n_50 & mul_74_11_n_30));
 assign n_1526 = ((n_1482 & ~n_1479) | (mul_74_11_n_37 & n_1479));
 assign n_1527 = (n_1484 ^ mul_74_11_n_42);
 assign n_1528 = ~(mul_74_11_n_38 ^ n_1286);
 assign n_1529 = ((n_1277 & ~mul_74_11_n_31) | (mul_74_11_n_41 & mul_74_11_n_31));
 assign n_1530 = ~((mul_74_11_n_49 & ~n_1286) | (n_1279 & n_1286));
 assign n_1531 = ((n_1484 & ~n_1280) | (mul_74_11_n_30 & n_1280));
 assign n_1532 = ~((mul_74_11_n_49 & ~n_1482) | (n_1279 & n_1482));
 assign n_1533 = ((n_1482 & ~n_1282) | (mul_74_11_n_37 & n_1282));
 assign n_1534 = ((n_1482 & ~n_1278) | (mul_74_11_n_37 & n_1278));
endmodule

