`timescale 1ps / 1ps
module dut_Mul2Add2Mul2u8u8u32Add2Mul2u29Add2u8u8Mul2u32Add2u8u8_4(
          in9,
          in8,
          in7,
          in6,
          in5,
          in4,
          in3,
          in2,
          in1,
          out1,
          clk
);
   input [7:0] in9;
   input [7:0] in8;
   input [31:0] in7;
   input [7:0] in6;
   input [7:0] in5;
   input [28:0] in4;
   input [31:0] in3;
   input [7:0] in2;
   input [7:0] in1;
   output [31:0] out1;
   input clk;
wire add_59_2_n_2, add_59_2_n_3, add_59_2_n_4, add_59_2_n_5, add_59_2_n_6,
     add_59_2_n_7, add_59_2_n_9, add_59_2_n_10, add_59_2_n_11, add_59_2_n_12,
     add_59_2_n_13, add_59_2_n_14, add_59_2_n_15, add_59_2_n_16, add_59_2_n_17,
     add_59_2_n_18, add_59_2_n_19, add_59_2_n_20, add_59_2_n_21, add_59_2_n_22,
     add_59_2_n_23, add_59_2_n_24, add_59_2_n_25, add_59_2_n_26, add_59_2_n_27,
     add_59_2_n_28, add_59_2_n_30, add_59_2_n_31, add_59_2_n_32, add_59_2_n_33,
     add_59_2_n_34, add_59_2_n_35, add_59_2_n_36, add_59_2_n_37, add_59_2_n_38,
     add_59_2_n_40, add_59_2_n_42, add_59_2_n_43, add_59_2_n_50, add_59_2_n_52,
     add_59_2_n_55, add_59_2_n_56, add_59_2_n_58, add_59_2_n_59, add_59_2_n_60,
     add_59_2_n_63, add_59_2_n_64, add_59_2_n_68, add_63_2_n_2, add_63_2_n_3,
     add_63_2_n_4, add_63_2_n_5, add_63_2_n_6, add_63_2_n_7, add_63_2_n_9,
     add_63_2_n_10, add_63_2_n_11, add_63_2_n_12, add_63_2_n_13, add_63_2_n_14,
     add_63_2_n_15, add_63_2_n_16, add_63_2_n_17, add_63_2_n_18, add_63_2_n_19,
     add_63_2_n_20, add_63_2_n_21, add_63_2_n_22, add_63_2_n_23, add_63_2_n_24,
     add_63_2_n_25, add_63_2_n_26, add_63_2_n_27, add_63_2_n_28, add_63_2_n_30,
     add_63_2_n_31, add_63_2_n_32, add_63_2_n_33, add_63_2_n_34, add_63_2_n_35,
     add_63_2_n_36, add_63_2_n_37, add_63_2_n_38, add_63_2_n_40, add_63_2_n_42,
     add_63_2_n_43, add_63_2_n_50, add_63_2_n_52, add_63_2_n_55, add_63_2_n_56,
     add_63_2_n_58, add_63_2_n_59, add_63_2_n_60, add_63_2_n_63, add_63_2_n_64,
     add_63_2_n_68, csa_tree_add_55_2_groupi_n_0, csa_tree_add_55_2_groupi_n_1,
     csa_tree_add_55_2_groupi_n_2, csa_tree_add_55_2_groupi_n_3,
     csa_tree_add_55_2_groupi_n_4, csa_tree_add_55_2_groupi_n_5,
     csa_tree_add_55_2_groupi_n_6, csa_tree_add_55_2_groupi_n_7,
     csa_tree_add_55_2_groupi_n_8, csa_tree_add_55_2_groupi_n_9,
     csa_tree_add_55_2_groupi_n_10, csa_tree_add_55_2_groupi_n_11,
     csa_tree_add_55_2_groupi_n_12, csa_tree_add_55_2_groupi_n_13,
     csa_tree_add_55_2_groupi_n_14, csa_tree_add_55_2_groupi_n_15,
     csa_tree_add_55_2_groupi_n_16, csa_tree_add_55_2_groupi_n_17,
     csa_tree_add_55_2_groupi_n_18, csa_tree_add_55_2_groupi_n_19,
     csa_tree_add_55_2_groupi_n_20, csa_tree_add_55_2_groupi_n_21,
     csa_tree_add_55_2_groupi_n_22, csa_tree_add_55_2_groupi_n_23,
     csa_tree_add_55_2_groupi_n_24, csa_tree_add_55_2_groupi_n_25,
     csa_tree_add_55_2_groupi_n_26, csa_tree_add_55_2_groupi_n_27,
     csa_tree_add_55_2_groupi_n_28, csa_tree_add_55_2_groupi_n_29,
     csa_tree_add_55_2_groupi_n_30, csa_tree_add_55_2_groupi_n_31,
     csa_tree_add_55_2_groupi_n_32, csa_tree_add_55_2_groupi_n_33,
     csa_tree_add_55_2_groupi_n_34, csa_tree_add_55_2_groupi_n_35,
     csa_tree_add_55_2_groupi_n_36, csa_tree_add_55_2_groupi_n_37,
     csa_tree_add_55_2_groupi_n_38, csa_tree_add_55_2_groupi_n_39,
     csa_tree_add_55_2_groupi_n_40, csa_tree_add_55_2_groupi_n_41,
     csa_tree_add_55_2_groupi_n_42, csa_tree_add_55_2_groupi_n_43,
     csa_tree_add_55_2_groupi_n_44, csa_tree_add_55_2_groupi_n_45,
     csa_tree_add_55_2_groupi_n_46, csa_tree_add_55_2_groupi_n_47,
     csa_tree_add_55_2_groupi_n_48, csa_tree_add_55_2_groupi_n_49,
     csa_tree_add_55_2_groupi_n_50, csa_tree_add_55_2_groupi_n_51,
     csa_tree_add_55_2_groupi_n_52, csa_tree_add_55_2_groupi_n_53,
     csa_tree_add_55_2_groupi_n_54, csa_tree_add_55_2_groupi_n_55,
     csa_tree_add_55_2_groupi_n_56, csa_tree_add_55_2_groupi_n_57,
     csa_tree_add_55_2_groupi_n_58, csa_tree_add_55_2_groupi_n_59,
     csa_tree_add_55_2_groupi_n_60, csa_tree_add_55_2_groupi_n_61,
     csa_tree_add_55_2_groupi_n_62, csa_tree_add_55_2_groupi_n_63,
     csa_tree_add_55_2_groupi_n_64, csa_tree_add_55_2_groupi_n_65,
     csa_tree_add_55_2_groupi_n_66, csa_tree_add_55_2_groupi_n_67,
     csa_tree_add_55_2_groupi_n_68, csa_tree_add_55_2_groupi_n_69,
     csa_tree_add_55_2_groupi_n_70, csa_tree_add_55_2_groupi_n_71,
     csa_tree_add_55_2_groupi_n_72, csa_tree_add_55_2_groupi_n_73,
     csa_tree_add_55_2_groupi_n_74, csa_tree_add_55_2_groupi_n_75,
     csa_tree_add_55_2_groupi_n_76, csa_tree_add_55_2_groupi_n_77,
     csa_tree_add_55_2_groupi_n_80, csa_tree_add_55_2_groupi_n_81,
     csa_tree_add_55_2_groupi_n_82, csa_tree_add_55_2_groupi_n_83,
     csa_tree_add_55_2_groupi_n_84, csa_tree_add_55_2_groupi_n_85,
     csa_tree_add_55_2_groupi_n_86, csa_tree_add_55_2_groupi_n_87,
     csa_tree_add_55_2_groupi_n_88, csa_tree_add_55_2_groupi_n_89,
     csa_tree_add_55_2_groupi_n_90, csa_tree_add_55_2_groupi_n_91,
     csa_tree_add_55_2_groupi_n_92, csa_tree_add_55_2_groupi_n_93,
     csa_tree_add_55_2_groupi_n_94, csa_tree_add_55_2_groupi_n_95,
     csa_tree_add_55_2_groupi_n_96, csa_tree_add_55_2_groupi_n_97,
     csa_tree_add_55_2_groupi_n_98, csa_tree_add_55_2_groupi_n_99,
     csa_tree_add_55_2_groupi_n_100, csa_tree_add_55_2_groupi_n_101,
     csa_tree_add_55_2_groupi_n_102, csa_tree_add_55_2_groupi_n_103,
     csa_tree_add_55_2_groupi_n_104, csa_tree_add_55_2_groupi_n_105,
     csa_tree_add_55_2_groupi_n_106, csa_tree_add_55_2_groupi_n_107,
     csa_tree_add_55_2_groupi_n_108, csa_tree_add_55_2_groupi_n_109,
     csa_tree_add_55_2_groupi_n_110, csa_tree_add_55_2_groupi_n_111,
     csa_tree_add_55_2_groupi_n_112, csa_tree_add_55_2_groupi_n_113,
     csa_tree_add_55_2_groupi_n_114, csa_tree_add_55_2_groupi_n_115,
     csa_tree_add_55_2_groupi_n_116, csa_tree_add_55_2_groupi_n_117,
     csa_tree_add_55_2_groupi_n_118, csa_tree_add_55_2_groupi_n_119,
     csa_tree_add_55_2_groupi_n_120, csa_tree_add_55_2_groupi_n_121,
     csa_tree_add_55_2_groupi_n_122, csa_tree_add_55_2_groupi_n_123,
     csa_tree_add_55_2_groupi_n_124, csa_tree_add_55_2_groupi_n_125,
     csa_tree_add_55_2_groupi_n_128, csa_tree_add_55_2_groupi_n_129,
     csa_tree_add_55_2_groupi_n_130, csa_tree_add_55_2_groupi_n_131,
     csa_tree_add_55_2_groupi_n_132, csa_tree_add_55_2_groupi_n_133,
     csa_tree_add_55_2_groupi_n_134, csa_tree_add_55_2_groupi_n_135,
     csa_tree_add_55_2_groupi_n_136, csa_tree_add_55_2_groupi_n_137,
     csa_tree_add_55_2_groupi_n_138, csa_tree_add_55_2_groupi_n_139,
     csa_tree_add_55_2_groupi_n_140, csa_tree_add_55_2_groupi_n_141,
     csa_tree_add_55_2_groupi_n_142, csa_tree_add_55_2_groupi_n_143,
     csa_tree_add_55_2_groupi_n_144, csa_tree_add_55_2_groupi_n_145,
     csa_tree_add_55_2_groupi_n_146, csa_tree_add_55_2_groupi_n_147,
     csa_tree_add_55_2_groupi_n_148, csa_tree_add_55_2_groupi_n_149,
     csa_tree_add_55_2_groupi_n_150, csa_tree_add_55_2_groupi_n_151,
     csa_tree_add_55_2_groupi_n_154, csa_tree_add_55_2_groupi_n_155,
     csa_tree_add_55_2_groupi_n_156, csa_tree_add_55_2_groupi_n_157,
     csa_tree_add_55_2_groupi_n_158, csa_tree_add_55_2_groupi_n_159,
     csa_tree_add_55_2_groupi_n_160, csa_tree_add_55_2_groupi_n_161,
     csa_tree_add_55_2_groupi_n_162, csa_tree_add_55_2_groupi_n_163,
     csa_tree_add_55_2_groupi_n_164, csa_tree_add_55_2_groupi_n_165,
     csa_tree_add_55_2_groupi_n_168, csa_tree_add_55_2_groupi_n_169,
     csa_tree_add_55_2_groupi_n_170, csa_tree_add_55_2_groupi_n_171,
     csa_tree_add_55_2_groupi_n_172, csa_tree_add_55_2_groupi_n_173,
     csa_tree_add_55_2_groupi_n_174, csa_tree_add_55_2_groupi_n_175,
     csa_tree_add_55_2_groupi_n_178, csa_tree_add_55_2_groupi_n_179,
     csa_tree_add_55_2_groupi_n_180, csa_tree_add_55_2_groupi_n_181,
     csa_tree_add_55_2_groupi_n_184, csa_tree_add_55_2_groupi_n_185,
     csa_tree_add_55_2_groupi_n_186, csa_tree_add_55_2_groupi_n_187,
     csa_tree_add_55_2_groupi_n_207, csa_tree_add_55_2_groupi_n_208,
     csa_tree_add_55_2_groupi_n_210, csa_tree_add_55_2_groupi_n_212,
     csa_tree_add_55_2_groupi_n_214, csa_tree_add_55_2_groupi_n_216,
     csa_tree_add_55_2_groupi_n_218, csa_tree_add_55_2_groupi_n_220,
     csa_tree_add_55_2_groupi_n_222, csa_tree_add_55_2_groupi_n_224,
     csa_tree_add_55_2_groupi_n_226, csa_tree_add_55_2_groupi_n_228,
     csa_tree_add_69_2_groupi_n_0, csa_tree_add_69_2_groupi_n_6,
     csa_tree_add_69_2_groupi_n_9, csa_tree_add_69_2_groupi_n_10,
     csa_tree_add_69_2_groupi_n_11, csa_tree_add_69_2_groupi_n_12,
     csa_tree_add_69_2_groupi_n_13, csa_tree_add_69_2_groupi_n_14,
     csa_tree_add_69_2_groupi_n_15, csa_tree_add_69_2_groupi_n_16,
     csa_tree_add_69_2_groupi_n_17, csa_tree_add_69_2_groupi_n_18,
     csa_tree_add_69_2_groupi_n_19, csa_tree_add_69_2_groupi_n_20,
     csa_tree_add_69_2_groupi_n_21, csa_tree_add_69_2_groupi_n_22,
     csa_tree_add_69_2_groupi_n_23, csa_tree_add_69_2_groupi_n_24,
     csa_tree_add_69_2_groupi_n_26, csa_tree_add_69_2_groupi_n_27,
     csa_tree_add_69_2_groupi_n_28, csa_tree_add_69_2_groupi_n_29,
     csa_tree_add_69_2_groupi_n_31, csa_tree_add_69_2_groupi_n_32,
     csa_tree_add_69_2_groupi_n_33, csa_tree_add_69_2_groupi_n_36,
     csa_tree_add_69_2_groupi_n_37, csa_tree_add_69_2_groupi_n_38,
     csa_tree_add_69_2_groupi_n_39, csa_tree_add_69_2_groupi_n_40,
     csa_tree_add_69_2_groupi_n_41, csa_tree_add_69_2_groupi_n_42,
     csa_tree_add_69_2_groupi_n_43, csa_tree_add_69_2_groupi_n_44,
     csa_tree_add_69_2_groupi_n_45, csa_tree_add_69_2_groupi_n_46,
     csa_tree_add_69_2_groupi_n_48, csa_tree_add_69_2_groupi_n_50,
     csa_tree_add_69_2_groupi_n_51, csa_tree_add_69_2_groupi_n_52,
     csa_tree_add_69_2_groupi_n_53, csa_tree_add_69_2_groupi_n_54,
     csa_tree_add_69_2_groupi_n_56, csa_tree_add_69_2_groupi_n_58,
     csa_tree_add_69_2_groupi_n_64, csa_tree_add_69_2_groupi_n_65,
     csa_tree_add_69_2_groupi_n_66, csa_tree_add_69_2_groupi_n_67,
     csa_tree_add_69_2_groupi_n_68, csa_tree_add_69_2_groupi_n_69,
     csa_tree_add_69_2_groupi_n_70, csa_tree_add_69_2_groupi_n_71,
     csa_tree_add_69_2_groupi_n_72, csa_tree_add_69_2_groupi_n_73,
     csa_tree_add_69_2_groupi_n_74, csa_tree_add_69_2_groupi_n_75,
     csa_tree_add_69_2_groupi_n_76, csa_tree_add_69_2_groupi_n_77,
     csa_tree_add_69_2_groupi_n_78, csa_tree_add_69_2_groupi_n_79,
     csa_tree_add_69_2_groupi_n_80, csa_tree_add_69_2_groupi_n_82,
     csa_tree_add_69_2_groupi_n_83, csa_tree_add_69_2_groupi_n_84,
     csa_tree_add_69_2_groupi_n_85, csa_tree_add_69_2_groupi_n_86,
     csa_tree_add_69_2_groupi_n_87, csa_tree_add_69_2_groupi_n_88,
     csa_tree_add_69_2_groupi_n_89, csa_tree_add_69_2_groupi_n_90,
     csa_tree_add_69_2_groupi_n_92, csa_tree_add_69_2_groupi_n_93,
     csa_tree_add_69_2_groupi_n_94, csa_tree_add_69_2_groupi_n_95,
     csa_tree_add_69_2_groupi_n_96, csa_tree_add_69_2_groupi_n_97,
     csa_tree_add_69_2_groupi_n_99, csa_tree_add_69_2_groupi_n_100,
     csa_tree_add_69_2_groupi_n_101, csa_tree_add_69_2_groupi_n_102,
     csa_tree_add_69_2_groupi_n_103, csa_tree_add_69_2_groupi_n_104,
     csa_tree_add_69_2_groupi_n_105, csa_tree_add_69_2_groupi_n_106,
     csa_tree_add_69_2_groupi_n_107, csa_tree_add_69_2_groupi_n_108,
     csa_tree_add_69_2_groupi_n_109, csa_tree_add_69_2_groupi_n_110,
     csa_tree_add_69_2_groupi_n_111, csa_tree_add_69_2_groupi_n_112,
     csa_tree_add_69_2_groupi_n_113, csa_tree_add_69_2_groupi_n_114,
     csa_tree_add_69_2_groupi_n_115, csa_tree_add_69_2_groupi_n_116,
     csa_tree_add_69_2_groupi_n_117, csa_tree_add_69_2_groupi_n_118,
     csa_tree_add_69_2_groupi_n_119, csa_tree_add_69_2_groupi_n_120,
     csa_tree_add_69_2_groupi_n_121, csa_tree_add_69_2_groupi_n_122,
     csa_tree_add_69_2_groupi_n_123, csa_tree_add_69_2_groupi_n_124,
     csa_tree_add_69_2_groupi_n_125, csa_tree_add_69_2_groupi_n_126,
     csa_tree_add_69_2_groupi_n_127, csa_tree_add_69_2_groupi_n_128,
     csa_tree_add_69_2_groupi_n_129, csa_tree_add_69_2_groupi_n_130,
     csa_tree_add_69_2_groupi_n_131, csa_tree_add_69_2_groupi_n_133,
     csa_tree_add_69_2_groupi_n_134, csa_tree_add_69_2_groupi_n_136,
     csa_tree_add_69_2_groupi_n_137, csa_tree_add_69_2_groupi_n_138,
     csa_tree_add_69_2_groupi_n_139, csa_tree_add_69_2_groupi_n_140,
     csa_tree_add_69_2_groupi_n_141, csa_tree_add_69_2_groupi_n_142,
     csa_tree_add_69_2_groupi_n_143, csa_tree_add_69_2_groupi_n_144,
     csa_tree_add_69_2_groupi_n_145, csa_tree_add_69_2_groupi_n_146,
     csa_tree_add_69_2_groupi_n_147, csa_tree_add_69_2_groupi_n_148,
     csa_tree_add_69_2_groupi_n_149, csa_tree_add_69_2_groupi_n_150,
     csa_tree_add_69_2_groupi_n_151, csa_tree_add_69_2_groupi_n_152,
     csa_tree_add_69_2_groupi_n_153, csa_tree_add_69_2_groupi_n_154,
     csa_tree_add_69_2_groupi_n_155, csa_tree_add_69_2_groupi_n_156,
     csa_tree_add_69_2_groupi_n_157, csa_tree_add_69_2_groupi_n_158,
     csa_tree_add_69_2_groupi_n_159, csa_tree_add_69_2_groupi_n_160,
     csa_tree_add_69_2_groupi_n_161, csa_tree_add_69_2_groupi_n_162,
     csa_tree_add_69_2_groupi_n_163, csa_tree_add_69_2_groupi_n_165,
     csa_tree_add_69_2_groupi_n_166, csa_tree_add_69_2_groupi_n_167,
     csa_tree_add_69_2_groupi_n_172, csa_tree_add_69_2_groupi_n_182,
     csa_tree_add_69_2_groupi_n_206, csa_tree_add_69_2_groupi_n_226,
     csa_tree_add_69_2_groupi_n_227, csa_tree_add_69_2_groupi_n_228,
     csa_tree_add_69_2_groupi_n_229, csa_tree_add_69_2_groupi_n_254,
     csa_tree_add_69_2_groupi_n_255, csa_tree_add_69_2_groupi_n_256,
     csa_tree_add_69_2_groupi_n_258, csa_tree_add_69_2_groupi_n_262,
     csa_tree_add_69_2_groupi_n_266, csa_tree_add_69_2_groupi_n_268,
     csa_tree_add_69_2_groupi_n_269, csa_tree_add_69_2_groupi_n_270,
     csa_tree_add_69_2_groupi_n_272, csa_tree_add_69_2_groupi_n_275,
     csa_tree_add_69_2_groupi_n_276, csa_tree_add_69_2_groupi_n_277,
     csa_tree_add_69_2_groupi_n_278, csa_tree_add_69_2_groupi_n_279,
     csa_tree_add_69_2_groupi_n_280, csa_tree_add_69_2_groupi_n_281,
     csa_tree_add_69_2_groupi_n_283, csa_tree_add_69_2_groupi_n_284,
     csa_tree_add_69_2_groupi_n_285, csa_tree_add_69_2_groupi_n_287,
     csa_tree_add_69_2_groupi_n_288, csa_tree_add_69_2_groupi_n_290,
     csa_tree_add_69_2_groupi_n_291, csa_tree_add_69_2_groupi_n_292,
     csa_tree_add_69_2_groupi_n_294, csa_tree_add_69_2_groupi_n_295,
     csa_tree_add_69_2_groupi_n_296, csa_tree_add_69_2_groupi_n_297,
     csa_tree_add_69_2_groupi_n_300, csa_tree_add_69_2_groupi_n_301,
     csa_tree_add_69_2_groupi_n_302, csa_tree_add_69_2_groupi_n_303,
     csa_tree_add_69_2_groupi_n_304, csa_tree_add_69_2_groupi_n_305,
     csa_tree_add_69_2_groupi_n_306, csa_tree_add_69_2_groupi_n_307,
     csa_tree_add_69_2_groupi_n_308, csa_tree_add_69_2_groupi_n_309,
     csa_tree_add_69_2_groupi_n_310, csa_tree_add_69_2_groupi_n_312,
     csa_tree_add_69_2_groupi_n_313, csa_tree_add_69_2_groupi_n_315,
     csa_tree_add_69_2_groupi_n_316, csa_tree_add_69_2_groupi_n_317,
     csa_tree_add_69_2_groupi_n_318, csa_tree_add_69_2_groupi_n_319,
     csa_tree_add_69_2_groupi_n_321, csa_tree_add_69_2_groupi_n_322,
     csa_tree_add_69_2_groupi_n_323, csa_tree_add_69_2_groupi_n_324,
     csa_tree_add_69_2_groupi_n_325, csa_tree_add_69_2_groupi_n_326,
     csa_tree_add_69_2_groupi_n_328, csa_tree_add_69_2_groupi_n_329,
     csa_tree_add_69_2_groupi_n_330, csa_tree_add_69_2_groupi_n_331,
     csa_tree_add_69_2_groupi_n_333, csa_tree_add_69_2_groupi_n_334,
     csa_tree_add_69_2_groupi_n_335, csa_tree_add_69_2_groupi_n_337,
     csa_tree_add_69_2_groupi_n_339, csa_tree_add_69_2_groupi_n_340,
     csa_tree_add_69_2_groupi_n_341, csa_tree_add_69_2_groupi_n_343,
     csa_tree_add_69_2_groupi_n_344, csa_tree_add_69_2_groupi_n_345,
     csa_tree_add_69_2_groupi_n_346, csa_tree_add_69_2_groupi_n_347,
     csa_tree_add_69_2_groupi_n_348, csa_tree_add_69_2_groupi_n_349,
     csa_tree_add_69_2_groupi_n_350, csa_tree_add_69_2_groupi_n_353,
     csa_tree_add_69_2_groupi_n_354, csa_tree_add_69_2_groupi_n_355,
     csa_tree_add_69_2_groupi_n_356, csa_tree_add_69_2_groupi_n_357,
     csa_tree_add_69_2_groupi_n_358, csa_tree_add_69_2_groupi_n_359,
     csa_tree_add_69_2_groupi_n_362, csa_tree_add_69_2_groupi_n_363,
     csa_tree_add_69_2_groupi_n_364, csa_tree_add_69_2_groupi_n_365,
     csa_tree_add_69_2_groupi_n_366, csa_tree_add_69_2_groupi_n_368,
     csa_tree_add_69_2_groupi_n_369, csa_tree_add_69_2_groupi_n_370,
     csa_tree_add_69_2_groupi_n_371, csa_tree_add_69_2_groupi_n_372,
     csa_tree_add_69_2_groupi_n_373, csa_tree_add_69_2_groupi_n_374,
     csa_tree_add_69_2_groupi_n_375, csa_tree_add_69_2_groupi_n_376,
     csa_tree_add_69_2_groupi_n_377, csa_tree_add_69_2_groupi_n_378,
     csa_tree_add_69_2_groupi_n_379, csa_tree_add_69_2_groupi_n_380,
     csa_tree_add_69_2_groupi_n_381, csa_tree_add_69_2_groupi_n_382,
     csa_tree_add_69_2_groupi_n_383, csa_tree_add_69_2_groupi_n_385,
     csa_tree_add_69_2_groupi_n_387, csa_tree_add_69_2_groupi_n_388,
     csa_tree_add_69_2_groupi_n_390, csa_tree_add_69_2_groupi_n_391,
     csa_tree_add_69_2_groupi_n_392, csa_tree_add_69_2_groupi_n_393,
     csa_tree_add_69_2_groupi_n_394, csa_tree_add_69_2_groupi_n_396,
     csa_tree_add_69_2_groupi_n_397, csa_tree_add_69_2_groupi_n_398,
     csa_tree_add_69_2_groupi_n_400, csa_tree_add_69_2_groupi_n_401,
     csa_tree_add_69_2_groupi_n_404, csa_tree_add_69_2_groupi_n_405,
     csa_tree_add_69_2_groupi_n_407, csa_tree_add_69_2_groupi_n_408,
     csa_tree_add_69_2_groupi_n_409, csa_tree_add_69_2_groupi_n_410,
     csa_tree_add_69_2_groupi_n_411, csa_tree_add_69_2_groupi_n_412,
     csa_tree_add_69_2_groupi_n_413, csa_tree_add_69_2_groupi_n_414,
     csa_tree_add_69_2_groupi_n_415, csa_tree_add_69_2_groupi_n_416,
     csa_tree_add_69_2_groupi_n_419, csa_tree_add_69_2_groupi_n_420,
     csa_tree_add_69_2_groupi_n_421, csa_tree_add_69_2_groupi_n_422,
     csa_tree_add_69_2_groupi_n_425, csa_tree_add_69_2_groupi_n_427,
     csa_tree_add_69_2_groupi_n_430, csa_tree_add_69_2_groupi_n_431,
     csa_tree_add_69_2_groupi_n_432, csa_tree_add_69_2_groupi_n_433,
     csa_tree_add_69_2_groupi_n_435, csa_tree_add_69_2_groupi_n_436,
     csa_tree_add_69_2_groupi_n_437, csa_tree_add_69_2_groupi_n_439,
     csa_tree_add_69_2_groupi_n_440, csa_tree_add_69_2_groupi_n_441,
     csa_tree_add_69_2_groupi_n_443, csa_tree_add_69_2_groupi_n_445,
     csa_tree_add_69_2_groupi_n_446, csa_tree_add_69_2_groupi_n_447,
     csa_tree_add_69_2_groupi_n_450, csa_tree_add_69_2_groupi_n_451,
     csa_tree_add_69_2_groupi_n_452, csa_tree_add_69_2_groupi_n_454,
     csa_tree_add_69_2_groupi_n_455, csa_tree_add_69_2_groupi_n_458,
     csa_tree_add_69_2_groupi_n_459, csa_tree_add_69_2_groupi_n_460,
     csa_tree_add_69_2_groupi_n_461, csa_tree_add_69_2_groupi_n_462,
     csa_tree_add_69_2_groupi_n_465, csa_tree_add_69_2_groupi_n_466,
     csa_tree_add_69_2_groupi_n_468, csa_tree_add_69_2_groupi_n_470,
     csa_tree_add_69_2_groupi_n_471, csa_tree_add_69_2_groupi_n_473,
     csa_tree_add_69_2_groupi_n_474, csa_tree_add_69_2_groupi_n_476,
     csa_tree_add_69_2_groupi_n_477, csa_tree_add_69_2_groupi_n_478,
     csa_tree_add_69_2_groupi_n_481, csa_tree_add_69_2_groupi_n_483,
     csa_tree_add_69_2_groupi_n_486, csa_tree_add_69_2_groupi_n_488,
     csa_tree_add_69_2_groupi_n_489, csa_tree_add_69_2_groupi_n_490,
     csa_tree_add_69_2_groupi_n_491, csa_tree_add_69_2_groupi_n_492,
     csa_tree_add_69_2_groupi_n_493, csa_tree_add_69_2_groupi_n_494,
     csa_tree_add_69_2_groupi_n_495, csa_tree_add_69_2_groupi_n_496,
     csa_tree_add_69_2_groupi_n_497, csa_tree_add_69_2_groupi_n_498,
     csa_tree_add_69_2_groupi_n_499, csa_tree_add_69_2_groupi_n_500,
     csa_tree_add_69_2_groupi_n_501, csa_tree_add_69_2_groupi_n_502,
     csa_tree_add_69_2_groupi_n_503, csa_tree_add_69_2_groupi_n_504,
     csa_tree_add_69_2_groupi_n_505, csa_tree_add_69_2_groupi_n_506,
     csa_tree_add_69_2_groupi_n_507, csa_tree_add_69_2_groupi_n_508,
     csa_tree_add_69_2_groupi_n_509, csa_tree_add_69_2_groupi_n_510,
     csa_tree_add_69_2_groupi_n_511, csa_tree_add_69_2_groupi_n_512,
     csa_tree_add_69_2_groupi_n_513, csa_tree_add_69_2_groupi_n_514,
     csa_tree_add_69_2_groupi_n_515, csa_tree_add_69_2_groupi_n_516,
     csa_tree_add_69_2_groupi_n_517, csa_tree_add_69_2_groupi_n_518,
     csa_tree_add_69_2_groupi_n_519, csa_tree_add_69_2_groupi_n_522,
     csa_tree_add_69_2_groupi_n_523, csa_tree_add_69_2_groupi_n_524,
     csa_tree_add_69_2_groupi_n_525, csa_tree_add_69_2_groupi_n_526,
     csa_tree_add_69_2_groupi_n_527, csa_tree_add_69_2_groupi_n_529,
     csa_tree_add_69_2_groupi_n_530, csa_tree_add_69_2_groupi_n_531,
     csa_tree_add_69_2_groupi_n_532, csa_tree_add_69_2_groupi_n_533,
     csa_tree_add_69_2_groupi_n_534, csa_tree_add_69_2_groupi_n_535,
     csa_tree_add_69_2_groupi_n_536, csa_tree_add_69_2_groupi_n_537,
     csa_tree_add_69_2_groupi_n_538, csa_tree_add_69_2_groupi_n_540,
     csa_tree_add_69_2_groupi_n_541, csa_tree_add_69_2_groupi_n_542,
     csa_tree_add_69_2_groupi_n_543, csa_tree_add_69_2_groupi_n_544,
     csa_tree_add_69_2_groupi_n_545, csa_tree_add_69_2_groupi_n_546,
     csa_tree_add_69_2_groupi_n_547, csa_tree_add_69_2_groupi_n_548,
     csa_tree_add_69_2_groupi_n_549, csa_tree_add_69_2_groupi_n_550,
     csa_tree_add_69_2_groupi_n_551, csa_tree_add_69_2_groupi_n_552,
     csa_tree_add_69_2_groupi_n_553, csa_tree_add_69_2_groupi_n_554,
     csa_tree_add_69_2_groupi_n_555, csa_tree_add_69_2_groupi_n_556,
     csa_tree_add_69_2_groupi_n_557, csa_tree_add_69_2_groupi_n_558,
     csa_tree_add_69_2_groupi_n_559, csa_tree_add_69_2_groupi_n_560,
     csa_tree_add_69_2_groupi_n_561, csa_tree_add_69_2_groupi_n_562,
     csa_tree_add_69_2_groupi_n_563, csa_tree_add_69_2_groupi_n_564,
     csa_tree_add_69_2_groupi_n_565, csa_tree_add_69_2_groupi_n_566,
     csa_tree_add_69_2_groupi_n_567, csa_tree_add_69_2_groupi_n_568,
     csa_tree_add_69_2_groupi_n_569, csa_tree_add_69_2_groupi_n_570,
     csa_tree_add_69_2_groupi_n_571, csa_tree_add_69_2_groupi_n_572,
     csa_tree_add_69_2_groupi_n_573, csa_tree_add_69_2_groupi_n_574,
     csa_tree_add_69_2_groupi_n_575, csa_tree_add_69_2_groupi_n_576,
     csa_tree_add_69_2_groupi_n_577, csa_tree_add_69_2_groupi_n_578,
     csa_tree_add_69_2_groupi_n_579, csa_tree_add_69_2_groupi_n_580,
     csa_tree_add_69_2_groupi_n_581, csa_tree_add_69_2_groupi_n_582,
     csa_tree_add_69_2_groupi_n_583, csa_tree_add_69_2_groupi_n_584,
     csa_tree_add_69_2_groupi_n_585, csa_tree_add_69_2_groupi_n_586,
     csa_tree_add_69_2_groupi_n_587, csa_tree_add_69_2_groupi_n_588,
     csa_tree_add_69_2_groupi_n_589, csa_tree_add_69_2_groupi_n_590,
     csa_tree_add_69_2_groupi_n_591, csa_tree_add_69_2_groupi_n_592,
     csa_tree_add_69_2_groupi_n_593, csa_tree_add_69_2_groupi_n_594,
     csa_tree_add_69_2_groupi_n_595, csa_tree_add_69_2_groupi_n_596,
     csa_tree_add_69_2_groupi_n_597, csa_tree_add_69_2_groupi_n_598,
     csa_tree_add_69_2_groupi_n_599, csa_tree_add_69_2_groupi_n_600,
     csa_tree_add_69_2_groupi_n_601, csa_tree_add_69_2_groupi_n_602,
     csa_tree_add_69_2_groupi_n_603, csa_tree_add_69_2_groupi_n_604,
     csa_tree_add_69_2_groupi_n_605, csa_tree_add_69_2_groupi_n_606,
     csa_tree_add_69_2_groupi_n_607, csa_tree_add_69_2_groupi_n_608,
     csa_tree_add_69_2_groupi_n_609, csa_tree_add_69_2_groupi_n_610,
     csa_tree_add_69_2_groupi_n_611, csa_tree_add_69_2_groupi_n_612,
     csa_tree_add_69_2_groupi_n_613, csa_tree_add_69_2_groupi_n_614,
     csa_tree_add_69_2_groupi_n_615, csa_tree_add_69_2_groupi_n_616,
     csa_tree_add_69_2_groupi_n_617, csa_tree_add_69_2_groupi_n_618,
     csa_tree_add_69_2_groupi_n_619, csa_tree_add_69_2_groupi_n_620,
     csa_tree_add_69_2_groupi_n_621, csa_tree_add_69_2_groupi_n_622,
     csa_tree_add_69_2_groupi_n_623, csa_tree_add_69_2_groupi_n_624,
     csa_tree_add_69_2_groupi_n_625, csa_tree_add_69_2_groupi_n_626,
     csa_tree_add_69_2_groupi_n_627, csa_tree_add_69_2_groupi_n_628,
     csa_tree_add_69_2_groupi_n_629, csa_tree_add_69_2_groupi_n_630,
     csa_tree_add_69_2_groupi_n_631, csa_tree_add_69_2_groupi_n_632,
     csa_tree_add_69_2_groupi_n_633, csa_tree_add_69_2_groupi_n_634,
     csa_tree_add_69_2_groupi_n_635, csa_tree_add_69_2_groupi_n_636,
     csa_tree_add_69_2_groupi_n_637, csa_tree_add_69_2_groupi_n_638,
     csa_tree_add_69_2_groupi_n_639, csa_tree_add_69_2_groupi_n_641,
     csa_tree_add_69_2_groupi_n_642, csa_tree_add_69_2_groupi_n_643,
     csa_tree_add_69_2_groupi_n_644, csa_tree_add_69_2_groupi_n_645,
     csa_tree_add_69_2_groupi_n_646, csa_tree_add_69_2_groupi_n_647,
     csa_tree_add_69_2_groupi_n_649, csa_tree_add_69_2_groupi_n_650,
     csa_tree_add_69_2_groupi_n_651, csa_tree_add_69_2_groupi_n_652,
     csa_tree_add_69_2_groupi_n_653, csa_tree_add_69_2_groupi_n_654,
     csa_tree_add_69_2_groupi_n_655, csa_tree_add_69_2_groupi_n_656,
     csa_tree_add_69_2_groupi_n_657, csa_tree_add_69_2_groupi_n_658,
     csa_tree_add_69_2_groupi_n_659, csa_tree_add_69_2_groupi_n_660,
     csa_tree_add_69_2_groupi_n_661, csa_tree_add_69_2_groupi_n_662,
     csa_tree_add_69_2_groupi_n_663, csa_tree_add_69_2_groupi_n_664,
     csa_tree_add_69_2_groupi_n_665, csa_tree_add_69_2_groupi_n_666,
     csa_tree_add_69_2_groupi_n_667, csa_tree_add_69_2_groupi_n_668,
     csa_tree_add_69_2_groupi_n_669, csa_tree_add_69_2_groupi_n_670,
     csa_tree_add_69_2_groupi_n_671, csa_tree_add_69_2_groupi_n_672,
     csa_tree_add_69_2_groupi_n_673, csa_tree_add_69_2_groupi_n_674,
     csa_tree_add_69_2_groupi_n_675, csa_tree_add_69_2_groupi_n_676,
     csa_tree_add_69_2_groupi_n_677, csa_tree_add_69_2_groupi_n_678,
     csa_tree_add_69_2_groupi_n_679, csa_tree_add_69_2_groupi_n_680,
     csa_tree_add_69_2_groupi_n_681, csa_tree_add_69_2_groupi_n_682,
     csa_tree_add_69_2_groupi_n_683, csa_tree_add_69_2_groupi_n_684,
     csa_tree_add_69_2_groupi_n_685, csa_tree_add_69_2_groupi_n_686,
     csa_tree_add_69_2_groupi_n_687, csa_tree_add_69_2_groupi_n_688,
     csa_tree_add_69_2_groupi_n_689, csa_tree_add_69_2_groupi_n_690,
     csa_tree_add_69_2_groupi_n_691, csa_tree_add_69_2_groupi_n_692,
     csa_tree_add_69_2_groupi_n_693, csa_tree_add_69_2_groupi_n_694,
     csa_tree_add_69_2_groupi_n_695, csa_tree_add_69_2_groupi_n_696,
     csa_tree_add_69_2_groupi_n_697, csa_tree_add_69_2_groupi_n_698,
     csa_tree_add_69_2_groupi_n_699, csa_tree_add_69_2_groupi_n_700,
     csa_tree_add_69_2_groupi_n_701, csa_tree_add_69_2_groupi_n_702,
     csa_tree_add_69_2_groupi_n_703, csa_tree_add_69_2_groupi_n_704,
     csa_tree_add_69_2_groupi_n_705, csa_tree_add_69_2_groupi_n_706,
     csa_tree_add_69_2_groupi_n_707, csa_tree_add_69_2_groupi_n_708,
     csa_tree_add_69_2_groupi_n_709, csa_tree_add_69_2_groupi_n_710,
     csa_tree_add_69_2_groupi_n_711, csa_tree_add_69_2_groupi_n_712,
     csa_tree_add_69_2_groupi_n_713, csa_tree_add_69_2_groupi_n_714,
     csa_tree_add_69_2_groupi_n_715, csa_tree_add_69_2_groupi_n_716,
     csa_tree_add_69_2_groupi_n_717, csa_tree_add_69_2_groupi_n_718,
     csa_tree_add_69_2_groupi_n_719, csa_tree_add_69_2_groupi_n_720,
     csa_tree_add_69_2_groupi_n_721, csa_tree_add_69_2_groupi_n_722,
     csa_tree_add_69_2_groupi_n_723, csa_tree_add_69_2_groupi_n_724,
     csa_tree_add_69_2_groupi_n_725, csa_tree_add_69_2_groupi_n_726,
     csa_tree_add_69_2_groupi_n_727, csa_tree_add_69_2_groupi_n_728,
     csa_tree_add_69_2_groupi_n_729, csa_tree_add_69_2_groupi_n_730,
     csa_tree_add_69_2_groupi_n_731, csa_tree_add_69_2_groupi_n_732,
     csa_tree_add_69_2_groupi_n_733, csa_tree_add_69_2_groupi_n_734,
     csa_tree_add_69_2_groupi_n_735, csa_tree_add_69_2_groupi_n_736,
     csa_tree_add_69_2_groupi_n_737, csa_tree_add_69_2_groupi_n_738,
     csa_tree_add_69_2_groupi_n_739, csa_tree_add_69_2_groupi_n_740,
     csa_tree_add_69_2_groupi_n_741, csa_tree_add_69_2_groupi_n_742,
     csa_tree_add_69_2_groupi_n_743, csa_tree_add_69_2_groupi_n_744,
     csa_tree_add_69_2_groupi_n_745, csa_tree_add_69_2_groupi_n_746,
     csa_tree_add_69_2_groupi_n_747, csa_tree_add_69_2_groupi_n_748,
     csa_tree_add_69_2_groupi_n_749, csa_tree_add_69_2_groupi_n_750,
     csa_tree_add_69_2_groupi_n_752, csa_tree_add_69_2_groupi_n_753,
     csa_tree_add_69_2_groupi_n_754, csa_tree_add_69_2_groupi_n_755,
     csa_tree_add_69_2_groupi_n_756, csa_tree_add_69_2_groupi_n_757,
     csa_tree_add_69_2_groupi_n_758, csa_tree_add_69_2_groupi_n_759,
     csa_tree_add_69_2_groupi_n_760, csa_tree_add_69_2_groupi_n_761,
     csa_tree_add_69_2_groupi_n_762, csa_tree_add_69_2_groupi_n_763,
     csa_tree_add_69_2_groupi_n_764, csa_tree_add_69_2_groupi_n_765,
     csa_tree_add_69_2_groupi_n_766, csa_tree_add_69_2_groupi_n_767,
     csa_tree_add_69_2_groupi_n_768, csa_tree_add_69_2_groupi_n_769,
     csa_tree_add_69_2_groupi_n_770, csa_tree_add_69_2_groupi_n_771,
     csa_tree_add_69_2_groupi_n_772, csa_tree_add_69_2_groupi_n_773,
     csa_tree_add_69_2_groupi_n_774, csa_tree_add_69_2_groupi_n_775,
     csa_tree_add_69_2_groupi_n_776, csa_tree_add_69_2_groupi_n_777,
     csa_tree_add_69_2_groupi_n_778, csa_tree_add_69_2_groupi_n_779,
     csa_tree_add_69_2_groupi_n_780, csa_tree_add_69_2_groupi_n_781,
     csa_tree_add_69_2_groupi_n_782, csa_tree_add_69_2_groupi_n_783,
     csa_tree_add_69_2_groupi_n_784, csa_tree_add_69_2_groupi_n_785,
     csa_tree_add_69_2_groupi_n_786, csa_tree_add_69_2_groupi_n_787,
     csa_tree_add_69_2_groupi_n_788, csa_tree_add_69_2_groupi_n_789,
     csa_tree_add_69_2_groupi_n_790, csa_tree_add_69_2_groupi_n_791,
     csa_tree_add_69_2_groupi_n_792, csa_tree_add_69_2_groupi_n_793,
     csa_tree_add_69_2_groupi_n_794, csa_tree_add_69_2_groupi_n_795,
     csa_tree_add_69_2_groupi_n_796, csa_tree_add_69_2_groupi_n_797,
     csa_tree_add_69_2_groupi_n_798, csa_tree_add_69_2_groupi_n_799,
     csa_tree_add_69_2_groupi_n_800, csa_tree_add_69_2_groupi_n_801,
     csa_tree_add_69_2_groupi_n_802, csa_tree_add_69_2_groupi_n_803,
     csa_tree_add_69_2_groupi_n_804, csa_tree_add_69_2_groupi_n_805,
     csa_tree_add_69_2_groupi_n_806, csa_tree_add_69_2_groupi_n_807,
     csa_tree_add_69_2_groupi_n_808, csa_tree_add_69_2_groupi_n_809,
     csa_tree_add_69_2_groupi_n_810, csa_tree_add_69_2_groupi_n_811,
     csa_tree_add_69_2_groupi_n_812, csa_tree_add_69_2_groupi_n_813,
     csa_tree_add_69_2_groupi_n_814, csa_tree_add_69_2_groupi_n_815,
     csa_tree_add_69_2_groupi_n_816, csa_tree_add_69_2_groupi_n_817,
     csa_tree_add_69_2_groupi_n_818, csa_tree_add_69_2_groupi_n_819,
     csa_tree_add_69_2_groupi_n_820, csa_tree_add_69_2_groupi_n_821,
     csa_tree_add_69_2_groupi_n_822, csa_tree_add_69_2_groupi_n_823,
     csa_tree_add_69_2_groupi_n_824, csa_tree_add_69_2_groupi_n_825,
     csa_tree_add_69_2_groupi_n_826, csa_tree_add_69_2_groupi_n_827,
     csa_tree_add_69_2_groupi_n_828, csa_tree_add_69_2_groupi_n_829,
     csa_tree_add_69_2_groupi_n_830, csa_tree_add_69_2_groupi_n_831,
     csa_tree_add_69_2_groupi_n_832, csa_tree_add_69_2_groupi_n_833,
     csa_tree_add_69_2_groupi_n_834, csa_tree_add_69_2_groupi_n_835,
     csa_tree_add_69_2_groupi_n_836, csa_tree_add_69_2_groupi_n_837,
     csa_tree_add_69_2_groupi_n_838, csa_tree_add_69_2_groupi_n_839,
     csa_tree_add_69_2_groupi_n_840, csa_tree_add_69_2_groupi_n_841,
     csa_tree_add_69_2_groupi_n_842, csa_tree_add_69_2_groupi_n_843,
     csa_tree_add_69_2_groupi_n_844, csa_tree_add_69_2_groupi_n_845,
     csa_tree_add_69_2_groupi_n_846, csa_tree_add_69_2_groupi_n_847,
     csa_tree_add_69_2_groupi_n_848, csa_tree_add_69_2_groupi_n_849,
     csa_tree_add_69_2_groupi_n_850, csa_tree_add_69_2_groupi_n_851,
     csa_tree_add_69_2_groupi_n_852, csa_tree_add_69_2_groupi_n_853,
     csa_tree_add_69_2_groupi_n_854, csa_tree_add_69_2_groupi_n_855,
     csa_tree_add_69_2_groupi_n_856, csa_tree_add_69_2_groupi_n_857,
     csa_tree_add_69_2_groupi_n_858, csa_tree_add_69_2_groupi_n_859,
     csa_tree_add_69_2_groupi_n_860, csa_tree_add_69_2_groupi_n_861,
     csa_tree_add_69_2_groupi_n_862, csa_tree_add_69_2_groupi_n_863,
     csa_tree_add_69_2_groupi_n_864, csa_tree_add_69_2_groupi_n_865,
     csa_tree_add_69_2_groupi_n_866, csa_tree_add_69_2_groupi_n_867,
     csa_tree_add_69_2_groupi_n_868, csa_tree_add_69_2_groupi_n_869,
     csa_tree_add_69_2_groupi_n_870, csa_tree_add_69_2_groupi_n_871,
     csa_tree_add_69_2_groupi_n_872, csa_tree_add_69_2_groupi_n_873,
     csa_tree_add_69_2_groupi_n_874, csa_tree_add_69_2_groupi_n_875,
     csa_tree_add_69_2_groupi_n_876, csa_tree_add_69_2_groupi_n_877,
     csa_tree_add_69_2_groupi_n_878, csa_tree_add_69_2_groupi_n_879,
     csa_tree_add_69_2_groupi_n_880, csa_tree_add_69_2_groupi_n_881,
     csa_tree_add_69_2_groupi_n_882, csa_tree_add_69_2_groupi_n_883,
     csa_tree_add_69_2_groupi_n_884, csa_tree_add_69_2_groupi_n_885,
     csa_tree_add_69_2_groupi_n_886, csa_tree_add_69_2_groupi_n_887,
     csa_tree_add_69_2_groupi_n_888, csa_tree_add_69_2_groupi_n_889,
     csa_tree_add_69_2_groupi_n_890, csa_tree_add_69_2_groupi_n_891,
     csa_tree_add_69_2_groupi_n_892, csa_tree_add_69_2_groupi_n_893,
     csa_tree_add_69_2_groupi_n_894, csa_tree_add_69_2_groupi_n_895,
     csa_tree_add_69_2_groupi_n_896, csa_tree_add_69_2_groupi_n_897,
     csa_tree_add_69_2_groupi_n_898, csa_tree_add_69_2_groupi_n_899,
     csa_tree_add_69_2_groupi_n_900, csa_tree_add_69_2_groupi_n_901,
     csa_tree_add_69_2_groupi_n_902, csa_tree_add_69_2_groupi_n_903,
     csa_tree_add_69_2_groupi_n_904, csa_tree_add_69_2_groupi_n_905,
     csa_tree_add_69_2_groupi_n_906, csa_tree_add_69_2_groupi_n_907,
     csa_tree_add_69_2_groupi_n_908, csa_tree_add_69_2_groupi_n_909,
     csa_tree_add_69_2_groupi_n_910, csa_tree_add_69_2_groupi_n_911,
     csa_tree_add_69_2_groupi_n_912, csa_tree_add_69_2_groupi_n_913,
     csa_tree_add_69_2_groupi_n_914, csa_tree_add_69_2_groupi_n_915,
     csa_tree_add_69_2_groupi_n_916, csa_tree_add_69_2_groupi_n_917,
     csa_tree_add_69_2_groupi_n_918, csa_tree_add_69_2_groupi_n_919,
     csa_tree_add_69_2_groupi_n_920, csa_tree_add_69_2_groupi_n_921,
     csa_tree_add_69_2_groupi_n_922, csa_tree_add_69_2_groupi_n_923,
     csa_tree_add_69_2_groupi_n_924, csa_tree_add_69_2_groupi_n_925,
     csa_tree_add_69_2_groupi_n_926, csa_tree_add_69_2_groupi_n_927,
     csa_tree_add_69_2_groupi_n_928, csa_tree_add_69_2_groupi_n_929,
     csa_tree_add_69_2_groupi_n_930, csa_tree_add_69_2_groupi_n_931,
     csa_tree_add_69_2_groupi_n_932, csa_tree_add_69_2_groupi_n_933,
     csa_tree_add_69_2_groupi_n_934, csa_tree_add_69_2_groupi_n_935,
     csa_tree_add_69_2_groupi_n_936, csa_tree_add_69_2_groupi_n_937,
     csa_tree_add_69_2_groupi_n_938, csa_tree_add_69_2_groupi_n_939,
     csa_tree_add_69_2_groupi_n_940, csa_tree_add_69_2_groupi_n_941,
     csa_tree_add_69_2_groupi_n_942, csa_tree_add_69_2_groupi_n_943,
     csa_tree_add_69_2_groupi_n_944, csa_tree_add_69_2_groupi_n_945,
     csa_tree_add_69_2_groupi_n_946, csa_tree_add_69_2_groupi_n_947,
     csa_tree_add_69_2_groupi_n_948, csa_tree_add_69_2_groupi_n_949,
     csa_tree_add_69_2_groupi_n_950, csa_tree_add_69_2_groupi_n_951,
     csa_tree_add_69_2_groupi_n_952, csa_tree_add_69_2_groupi_n_953,
     csa_tree_add_69_2_groupi_n_954, csa_tree_add_69_2_groupi_n_955,
     csa_tree_add_69_2_groupi_n_956, csa_tree_add_69_2_groupi_n_957,
     csa_tree_add_69_2_groupi_n_958, csa_tree_add_69_2_groupi_n_959,
     csa_tree_add_69_2_groupi_n_960, csa_tree_add_69_2_groupi_n_961,
     csa_tree_add_69_2_groupi_n_962, csa_tree_add_69_2_groupi_n_963,
     csa_tree_add_69_2_groupi_n_964, csa_tree_add_69_2_groupi_n_965,
     csa_tree_add_69_2_groupi_n_966, csa_tree_add_69_2_groupi_n_967,
     csa_tree_add_69_2_groupi_n_968, csa_tree_add_69_2_groupi_n_969,
     csa_tree_add_69_2_groupi_n_970, csa_tree_add_69_2_groupi_n_971,
     csa_tree_add_69_2_groupi_n_972, csa_tree_add_69_2_groupi_n_973,
     csa_tree_add_69_2_groupi_n_974, csa_tree_add_69_2_groupi_n_975,
     csa_tree_add_69_2_groupi_n_976, csa_tree_add_69_2_groupi_n_977,
     csa_tree_add_69_2_groupi_n_978, csa_tree_add_69_2_groupi_n_979,
     csa_tree_add_69_2_groupi_n_980, csa_tree_add_69_2_groupi_n_981,
     csa_tree_add_69_2_groupi_n_982, csa_tree_add_69_2_groupi_n_983,
     csa_tree_add_69_2_groupi_n_984, csa_tree_add_69_2_groupi_n_985,
     csa_tree_add_69_2_groupi_n_987, csa_tree_add_69_2_groupi_n_988,
     csa_tree_add_69_2_groupi_n_989, csa_tree_add_69_2_groupi_n_990,
     csa_tree_add_69_2_groupi_n_991, csa_tree_add_69_2_groupi_n_992,
     csa_tree_add_69_2_groupi_n_993, csa_tree_add_69_2_groupi_n_994,
     csa_tree_add_69_2_groupi_n_995, csa_tree_add_69_2_groupi_n_997,
     csa_tree_add_69_2_groupi_n_998, csa_tree_add_69_2_groupi_n_999,
     csa_tree_add_69_2_groupi_n_1000, csa_tree_add_69_2_groupi_n_1001,
     csa_tree_add_69_2_groupi_n_1003, csa_tree_add_69_2_groupi_n_1004,
     csa_tree_add_69_2_groupi_n_1005, csa_tree_add_69_2_groupi_n_1007,
     csa_tree_add_69_2_groupi_n_1008, csa_tree_add_69_2_groupi_n_1009,
     csa_tree_add_69_2_groupi_n_1010, csa_tree_add_69_2_groupi_n_1011,
     csa_tree_add_69_2_groupi_n_1012, csa_tree_add_69_2_groupi_n_1013,
     csa_tree_add_69_2_groupi_n_1015, csa_tree_add_69_2_groupi_n_1016,
     csa_tree_add_69_2_groupi_n_1017, csa_tree_add_69_2_groupi_n_1018,
     csa_tree_add_69_2_groupi_n_1019, csa_tree_add_69_2_groupi_n_1020,
     csa_tree_add_69_2_groupi_n_1021, csa_tree_add_69_2_groupi_n_1023,
     csa_tree_add_69_2_groupi_n_1024, csa_tree_add_69_2_groupi_n_1025,
     csa_tree_add_69_2_groupi_n_1027, csa_tree_add_69_2_groupi_n_1028,
     csa_tree_add_69_2_groupi_n_1029, csa_tree_add_69_2_groupi_n_1030,
     csa_tree_add_69_2_groupi_n_1031, csa_tree_add_69_2_groupi_n_1032,
     csa_tree_add_69_2_groupi_n_1033, csa_tree_add_69_2_groupi_n_1034,
     csa_tree_add_69_2_groupi_n_1035, csa_tree_add_69_2_groupi_n_1036,
     csa_tree_add_69_2_groupi_n_1037, csa_tree_add_69_2_groupi_n_1038,
     csa_tree_add_69_2_groupi_n_1039, csa_tree_add_69_2_groupi_n_1040,
     csa_tree_add_69_2_groupi_n_1041, csa_tree_add_69_2_groupi_n_1042,
     csa_tree_add_69_2_groupi_n_1043, csa_tree_add_69_2_groupi_n_1044,
     csa_tree_add_69_2_groupi_n_1045, csa_tree_add_69_2_groupi_n_1046,
     csa_tree_add_69_2_groupi_n_1047, csa_tree_add_69_2_groupi_n_1048,
     csa_tree_add_69_2_groupi_n_1049, csa_tree_add_69_2_groupi_n_1050,
     csa_tree_add_69_2_groupi_n_1051, csa_tree_add_69_2_groupi_n_1052,
     csa_tree_add_69_2_groupi_n_1053, csa_tree_add_69_2_groupi_n_1054,
     csa_tree_add_69_2_groupi_n_1055, csa_tree_add_69_2_groupi_n_1056,
     csa_tree_add_69_2_groupi_n_1057, csa_tree_add_69_2_groupi_n_1058,
     csa_tree_add_69_2_groupi_n_1059, csa_tree_add_69_2_groupi_n_1060,
     csa_tree_add_69_2_groupi_n_1061, csa_tree_add_69_2_groupi_n_1062,
     csa_tree_add_69_2_groupi_n_1063, csa_tree_add_69_2_groupi_n_1064,
     csa_tree_add_69_2_groupi_n_1065, csa_tree_add_69_2_groupi_n_1066,
     csa_tree_add_69_2_groupi_n_1067, csa_tree_add_69_2_groupi_n_1068,
     csa_tree_add_69_2_groupi_n_1069, csa_tree_add_69_2_groupi_n_1070,
     csa_tree_add_69_2_groupi_n_1071, csa_tree_add_69_2_groupi_n_1072,
     csa_tree_add_69_2_groupi_n_1073, csa_tree_add_69_2_groupi_n_1074,
     csa_tree_add_69_2_groupi_n_1075, csa_tree_add_69_2_groupi_n_1076,
     csa_tree_add_69_2_groupi_n_1077, csa_tree_add_69_2_groupi_n_1078,
     csa_tree_add_69_2_groupi_n_1079, csa_tree_add_69_2_groupi_n_1081,
     csa_tree_add_69_2_groupi_n_1082, csa_tree_add_69_2_groupi_n_1083,
     csa_tree_add_69_2_groupi_n_1084, csa_tree_add_69_2_groupi_n_1085,
     csa_tree_add_69_2_groupi_n_1086, csa_tree_add_69_2_groupi_n_1087,
     csa_tree_add_69_2_groupi_n_1088, csa_tree_add_69_2_groupi_n_1089,
     csa_tree_add_69_2_groupi_n_1090, csa_tree_add_69_2_groupi_n_1091,
     csa_tree_add_69_2_groupi_n_1092, csa_tree_add_69_2_groupi_n_1093,
     csa_tree_add_69_2_groupi_n_1094, csa_tree_add_69_2_groupi_n_1095,
     csa_tree_add_69_2_groupi_n_1096, csa_tree_add_69_2_groupi_n_1097,
     csa_tree_add_69_2_groupi_n_1098, csa_tree_add_69_2_groupi_n_1099,
     csa_tree_add_69_2_groupi_n_1100, csa_tree_add_69_2_groupi_n_1101,
     csa_tree_add_69_2_groupi_n_1102, csa_tree_add_69_2_groupi_n_1103,
     csa_tree_add_69_2_groupi_n_1104, csa_tree_add_69_2_groupi_n_1105,
     csa_tree_add_69_2_groupi_n_1106, csa_tree_add_69_2_groupi_n_1107,
     csa_tree_add_69_2_groupi_n_1108, csa_tree_add_69_2_groupi_n_1109,
     csa_tree_add_69_2_groupi_n_1110, csa_tree_add_69_2_groupi_n_1111,
     csa_tree_add_69_2_groupi_n_1112, csa_tree_add_69_2_groupi_n_1113,
     csa_tree_add_69_2_groupi_n_1114, csa_tree_add_69_2_groupi_n_1115,
     csa_tree_add_69_2_groupi_n_1116, csa_tree_add_69_2_groupi_n_1117,
     csa_tree_add_69_2_groupi_n_1118, csa_tree_add_69_2_groupi_n_1119,
     csa_tree_add_69_2_groupi_n_1120, csa_tree_add_69_2_groupi_n_1121,
     csa_tree_add_69_2_groupi_n_1122, csa_tree_add_69_2_groupi_n_1123,
     csa_tree_add_69_2_groupi_n_1124, csa_tree_add_69_2_groupi_n_1125,
     csa_tree_add_69_2_groupi_n_1126, csa_tree_add_69_2_groupi_n_1127,
     csa_tree_add_69_2_groupi_n_1128, csa_tree_add_69_2_groupi_n_1129,
     csa_tree_add_69_2_groupi_n_1130, csa_tree_add_69_2_groupi_n_1131,
     csa_tree_add_69_2_groupi_n_1132, csa_tree_add_69_2_groupi_n_1133,
     csa_tree_add_69_2_groupi_n_1134, csa_tree_add_69_2_groupi_n_1135,
     csa_tree_add_69_2_groupi_n_1136, csa_tree_add_69_2_groupi_n_1137,
     csa_tree_add_69_2_groupi_n_1138, csa_tree_add_69_2_groupi_n_1139,
     csa_tree_add_69_2_groupi_n_1140, csa_tree_add_69_2_groupi_n_1141,
     csa_tree_add_69_2_groupi_n_1142, csa_tree_add_69_2_groupi_n_1143,
     csa_tree_add_69_2_groupi_n_1144, csa_tree_add_69_2_groupi_n_1145,
     csa_tree_add_69_2_groupi_n_1146, csa_tree_add_69_2_groupi_n_1147,
     csa_tree_add_69_2_groupi_n_1148, csa_tree_add_69_2_groupi_n_1149,
     csa_tree_add_69_2_groupi_n_1150, csa_tree_add_69_2_groupi_n_1151,
     csa_tree_add_69_2_groupi_n_1152, csa_tree_add_69_2_groupi_n_1153,
     csa_tree_add_69_2_groupi_n_1154, csa_tree_add_69_2_groupi_n_1155,
     csa_tree_add_69_2_groupi_n_1156, csa_tree_add_69_2_groupi_n_1157,
     csa_tree_add_69_2_groupi_n_1158, csa_tree_add_69_2_groupi_n_1159,
     csa_tree_add_69_2_groupi_n_1160, csa_tree_add_69_2_groupi_n_1161,
     csa_tree_add_69_2_groupi_n_1162, csa_tree_add_69_2_groupi_n_1163,
     csa_tree_add_69_2_groupi_n_1164, csa_tree_add_69_2_groupi_n_1165,
     csa_tree_add_69_2_groupi_n_1166, csa_tree_add_69_2_groupi_n_1167,
     csa_tree_add_69_2_groupi_n_1168, csa_tree_add_69_2_groupi_n_1169,
     csa_tree_add_69_2_groupi_n_1170, csa_tree_add_69_2_groupi_n_1171,
     csa_tree_add_69_2_groupi_n_1172, csa_tree_add_69_2_groupi_n_1173,
     csa_tree_add_69_2_groupi_n_1174, csa_tree_add_69_2_groupi_n_1175,
     csa_tree_add_69_2_groupi_n_1176, csa_tree_add_69_2_groupi_n_1177,
     csa_tree_add_69_2_groupi_n_1178, csa_tree_add_69_2_groupi_n_1179,
     csa_tree_add_69_2_groupi_n_1180, csa_tree_add_69_2_groupi_n_1181,
     csa_tree_add_69_2_groupi_n_1182, csa_tree_add_69_2_groupi_n_1183,
     csa_tree_add_69_2_groupi_n_1184, csa_tree_add_69_2_groupi_n_1185,
     csa_tree_add_69_2_groupi_n_1186, csa_tree_add_69_2_groupi_n_1187,
     csa_tree_add_69_2_groupi_n_1188, csa_tree_add_69_2_groupi_n_1189,
     csa_tree_add_69_2_groupi_n_1190, csa_tree_add_69_2_groupi_n_1191,
     csa_tree_add_69_2_groupi_n_1192, csa_tree_add_69_2_groupi_n_1193,
     csa_tree_add_69_2_groupi_n_1194, csa_tree_add_69_2_groupi_n_1195,
     csa_tree_add_69_2_groupi_n_1196, csa_tree_add_69_2_groupi_n_1197,
     csa_tree_add_69_2_groupi_n_1198, csa_tree_add_69_2_groupi_n_1199,
     csa_tree_add_69_2_groupi_n_1200, csa_tree_add_69_2_groupi_n_1201,
     csa_tree_add_69_2_groupi_n_1202, csa_tree_add_69_2_groupi_n_1203,
     csa_tree_add_69_2_groupi_n_1205, csa_tree_add_69_2_groupi_n_1206,
     csa_tree_add_69_2_groupi_n_1207, csa_tree_add_69_2_groupi_n_1208,
     csa_tree_add_69_2_groupi_n_1209, csa_tree_add_69_2_groupi_n_1210,
     csa_tree_add_69_2_groupi_n_1211, csa_tree_add_69_2_groupi_n_1212,
     csa_tree_add_69_2_groupi_n_1213, csa_tree_add_69_2_groupi_n_1214,
     csa_tree_add_69_2_groupi_n_1215, csa_tree_add_69_2_groupi_n_1216,
     csa_tree_add_69_2_groupi_n_1217, csa_tree_add_69_2_groupi_n_1218,
     csa_tree_add_69_2_groupi_n_1219, csa_tree_add_69_2_groupi_n_1220,
     csa_tree_add_69_2_groupi_n_1221, csa_tree_add_69_2_groupi_n_1222,
     csa_tree_add_69_2_groupi_n_1223, csa_tree_add_69_2_groupi_n_1224,
     csa_tree_add_69_2_groupi_n_1225, csa_tree_add_69_2_groupi_n_1226,
     csa_tree_add_69_2_groupi_n_1227, csa_tree_add_69_2_groupi_n_1228,
     csa_tree_add_69_2_groupi_n_1229, csa_tree_add_69_2_groupi_n_1230,
     csa_tree_add_69_2_groupi_n_1231, csa_tree_add_69_2_groupi_n_1232,
     csa_tree_add_69_2_groupi_n_1233, csa_tree_add_69_2_groupi_n_1234,
     csa_tree_add_69_2_groupi_n_1235, csa_tree_add_69_2_groupi_n_1236,
     csa_tree_add_69_2_groupi_n_1237, csa_tree_add_69_2_groupi_n_1238,
     csa_tree_add_69_2_groupi_n_1239, csa_tree_add_69_2_groupi_n_1240,
     csa_tree_add_69_2_groupi_n_1241, csa_tree_add_69_2_groupi_n_1242,
     csa_tree_add_69_2_groupi_n_1243, csa_tree_add_69_2_groupi_n_1244,
     csa_tree_add_69_2_groupi_n_1245, csa_tree_add_69_2_groupi_n_1246,
     csa_tree_add_69_2_groupi_n_1247, csa_tree_add_69_2_groupi_n_1248,
     csa_tree_add_69_2_groupi_n_1249, csa_tree_add_69_2_groupi_n_1250,
     csa_tree_add_69_2_groupi_n_1251, csa_tree_add_69_2_groupi_n_1252,
     csa_tree_add_69_2_groupi_n_1253, csa_tree_add_69_2_groupi_n_1254,
     csa_tree_add_69_2_groupi_n_1255, csa_tree_add_69_2_groupi_n_1256,
     csa_tree_add_69_2_groupi_n_1257, csa_tree_add_69_2_groupi_n_1258,
     csa_tree_add_69_2_groupi_n_1259, csa_tree_add_69_2_groupi_n_1260,
     csa_tree_add_69_2_groupi_n_1261, csa_tree_add_69_2_groupi_n_1262,
     csa_tree_add_69_2_groupi_n_1263, csa_tree_add_69_2_groupi_n_1264,
     csa_tree_add_69_2_groupi_n_1265, csa_tree_add_69_2_groupi_n_1266,
     csa_tree_add_69_2_groupi_n_1267, csa_tree_add_69_2_groupi_n_1268,
     csa_tree_add_69_2_groupi_n_1269, csa_tree_add_69_2_groupi_n_1270,
     csa_tree_add_69_2_groupi_n_1271, csa_tree_add_69_2_groupi_n_1272,
     csa_tree_add_69_2_groupi_n_1273, csa_tree_add_69_2_groupi_n_1274,
     csa_tree_add_69_2_groupi_n_1275, csa_tree_add_69_2_groupi_n_1276,
     csa_tree_add_69_2_groupi_n_1277, csa_tree_add_69_2_groupi_n_1278,
     csa_tree_add_69_2_groupi_n_1279, csa_tree_add_69_2_groupi_n_1280,
     csa_tree_add_69_2_groupi_n_1281, csa_tree_add_69_2_groupi_n_1282,
     csa_tree_add_69_2_groupi_n_1283, csa_tree_add_69_2_groupi_n_1284,
     csa_tree_add_69_2_groupi_n_1285, csa_tree_add_69_2_groupi_n_1286,
     csa_tree_add_69_2_groupi_n_1287, csa_tree_add_69_2_groupi_n_1288,
     csa_tree_add_69_2_groupi_n_1289, csa_tree_add_69_2_groupi_n_1290,
     csa_tree_add_69_2_groupi_n_1291, csa_tree_add_69_2_groupi_n_1292,
     csa_tree_add_69_2_groupi_n_1293, csa_tree_add_69_2_groupi_n_1294,
     csa_tree_add_69_2_groupi_n_1297, csa_tree_add_69_2_groupi_n_1298,
     csa_tree_add_69_2_groupi_n_1299, csa_tree_add_69_2_groupi_n_1300,
     csa_tree_add_69_2_groupi_n_1301, csa_tree_add_69_2_groupi_n_1303,
     csa_tree_add_69_2_groupi_n_1304, csa_tree_add_69_2_groupi_n_1305,
     csa_tree_add_69_2_groupi_n_1306, csa_tree_add_69_2_groupi_n_1307,
     csa_tree_add_69_2_groupi_n_1308, csa_tree_add_69_2_groupi_n_1309,
     csa_tree_add_69_2_groupi_n_1310, csa_tree_add_69_2_groupi_n_1311,
     csa_tree_add_69_2_groupi_n_1312, csa_tree_add_69_2_groupi_n_1313,
     csa_tree_add_69_2_groupi_n_1314, csa_tree_add_69_2_groupi_n_1315,
     csa_tree_add_69_2_groupi_n_1316, csa_tree_add_69_2_groupi_n_1317,
     csa_tree_add_69_2_groupi_n_1318, csa_tree_add_69_2_groupi_n_1319,
     csa_tree_add_69_2_groupi_n_1320, csa_tree_add_69_2_groupi_n_1321,
     csa_tree_add_69_2_groupi_n_1322, csa_tree_add_69_2_groupi_n_1323,
     csa_tree_add_69_2_groupi_n_1324, csa_tree_add_69_2_groupi_n_1325,
     csa_tree_add_69_2_groupi_n_1326, csa_tree_add_69_2_groupi_n_1327,
     csa_tree_add_69_2_groupi_n_1328, csa_tree_add_69_2_groupi_n_1329,
     csa_tree_add_69_2_groupi_n_1330, csa_tree_add_69_2_groupi_n_1331,
     csa_tree_add_69_2_groupi_n_1332, csa_tree_add_69_2_groupi_n_1333,
     csa_tree_add_69_2_groupi_n_1334, csa_tree_add_69_2_groupi_n_1335,
     csa_tree_add_69_2_groupi_n_1336, csa_tree_add_69_2_groupi_n_1337,
     csa_tree_add_69_2_groupi_n_1338, csa_tree_add_69_2_groupi_n_1339,
     csa_tree_add_69_2_groupi_n_1340, csa_tree_add_69_2_groupi_n_1341,
     csa_tree_add_69_2_groupi_n_1342, csa_tree_add_69_2_groupi_n_1343,
     csa_tree_add_69_2_groupi_n_1344, csa_tree_add_69_2_groupi_n_1345,
     csa_tree_add_69_2_groupi_n_1346, csa_tree_add_69_2_groupi_n_1347,
     csa_tree_add_69_2_groupi_n_1348, csa_tree_add_69_2_groupi_n_1349,
     csa_tree_add_69_2_groupi_n_1350, csa_tree_add_69_2_groupi_n_1351,
     csa_tree_add_69_2_groupi_n_1352, csa_tree_add_69_2_groupi_n_1353,
     csa_tree_add_69_2_groupi_n_1354, csa_tree_add_69_2_groupi_n_1355,
     csa_tree_add_69_2_groupi_n_1356, csa_tree_add_69_2_groupi_n_1357,
     csa_tree_add_69_2_groupi_n_1358, csa_tree_add_69_2_groupi_n_1359,
     csa_tree_add_69_2_groupi_n_1360, csa_tree_add_69_2_groupi_n_1361,
     csa_tree_add_69_2_groupi_n_1362, csa_tree_add_69_2_groupi_n_1363,
     csa_tree_add_69_2_groupi_n_1364, csa_tree_add_69_2_groupi_n_1365,
     csa_tree_add_69_2_groupi_n_1366, csa_tree_add_69_2_groupi_n_1367,
     csa_tree_add_69_2_groupi_n_1368, csa_tree_add_69_2_groupi_n_1369,
     csa_tree_add_69_2_groupi_n_1370, csa_tree_add_69_2_groupi_n_1371,
     csa_tree_add_69_2_groupi_n_1372, csa_tree_add_69_2_groupi_n_1373,
     csa_tree_add_69_2_groupi_n_1374, csa_tree_add_69_2_groupi_n_1375,
     csa_tree_add_69_2_groupi_n_1376, csa_tree_add_69_2_groupi_n_1377,
     csa_tree_add_69_2_groupi_n_1378, csa_tree_add_69_2_groupi_n_1379,
     csa_tree_add_69_2_groupi_n_1380, csa_tree_add_69_2_groupi_n_1381,
     csa_tree_add_69_2_groupi_n_1382, csa_tree_add_69_2_groupi_n_1383,
     csa_tree_add_69_2_groupi_n_1384, csa_tree_add_69_2_groupi_n_1385,
     csa_tree_add_69_2_groupi_n_1386, csa_tree_add_69_2_groupi_n_1387,
     csa_tree_add_69_2_groupi_n_1388, csa_tree_add_69_2_groupi_n_1389,
     csa_tree_add_69_2_groupi_n_1390, csa_tree_add_69_2_groupi_n_1391,
     csa_tree_add_69_2_groupi_n_1392, csa_tree_add_69_2_groupi_n_1393,
     csa_tree_add_69_2_groupi_n_1394, csa_tree_add_69_2_groupi_n_1395,
     csa_tree_add_69_2_groupi_n_1396, csa_tree_add_69_2_groupi_n_1397,
     csa_tree_add_69_2_groupi_n_1398, csa_tree_add_69_2_groupi_n_1399,
     csa_tree_add_69_2_groupi_n_1400, csa_tree_add_69_2_groupi_n_1401,
     csa_tree_add_69_2_groupi_n_1402, csa_tree_add_69_2_groupi_n_1403,
     csa_tree_add_69_2_groupi_n_1404, csa_tree_add_69_2_groupi_n_1405,
     csa_tree_add_69_2_groupi_n_1406, csa_tree_add_69_2_groupi_n_1407,
     csa_tree_add_69_2_groupi_n_1408, csa_tree_add_69_2_groupi_n_1409,
     csa_tree_add_69_2_groupi_n_1410, csa_tree_add_69_2_groupi_n_1411,
     csa_tree_add_69_2_groupi_n_1412, csa_tree_add_69_2_groupi_n_1413,
     csa_tree_add_69_2_groupi_n_1414, csa_tree_add_69_2_groupi_n_1417,
     csa_tree_add_69_2_groupi_n_1418, csa_tree_add_69_2_groupi_n_1420,
     csa_tree_add_69_2_groupi_n_1421, csa_tree_add_69_2_groupi_n_1424,
     csa_tree_add_69_2_groupi_n_1425, csa_tree_add_69_2_groupi_n_1427,
     csa_tree_add_69_2_groupi_n_1428, csa_tree_add_69_2_groupi_n_1429,
     csa_tree_add_69_2_groupi_n_1430, csa_tree_add_69_2_groupi_n_1431,
     csa_tree_add_69_2_groupi_n_1432, csa_tree_add_69_2_groupi_n_1433,
     csa_tree_add_69_2_groupi_n_1434, csa_tree_add_69_2_groupi_n_1435,
     csa_tree_add_69_2_groupi_n_1436, csa_tree_add_69_2_groupi_n_1437,
     csa_tree_add_69_2_groupi_n_1438, csa_tree_add_69_2_groupi_n_1439,
     csa_tree_add_69_2_groupi_n_1440, csa_tree_add_69_2_groupi_n_1441,
     csa_tree_add_69_2_groupi_n_1442, csa_tree_add_69_2_groupi_n_1443,
     csa_tree_add_69_2_groupi_n_1444, csa_tree_add_69_2_groupi_n_1445,
     csa_tree_add_69_2_groupi_n_1446, csa_tree_add_69_2_groupi_n_1447,
     csa_tree_add_69_2_groupi_n_1448, csa_tree_add_69_2_groupi_n_1449,
     csa_tree_add_69_2_groupi_n_1450, csa_tree_add_69_2_groupi_n_1451,
     csa_tree_add_69_2_groupi_n_1452, csa_tree_add_69_2_groupi_n_1453,
     csa_tree_add_69_2_groupi_n_1454, csa_tree_add_69_2_groupi_n_1455,
     csa_tree_add_69_2_groupi_n_1456, csa_tree_add_69_2_groupi_n_1457,
     csa_tree_add_69_2_groupi_n_1458, csa_tree_add_69_2_groupi_n_1459,
     csa_tree_add_69_2_groupi_n_1460, csa_tree_add_69_2_groupi_n_1461,
     csa_tree_add_69_2_groupi_n_1462, csa_tree_add_69_2_groupi_n_1463,
     csa_tree_add_69_2_groupi_n_1464, csa_tree_add_69_2_groupi_n_1466,
     csa_tree_add_69_2_groupi_n_1467, csa_tree_add_69_2_groupi_n_1468,
     csa_tree_add_69_2_groupi_n_1469, csa_tree_add_69_2_groupi_n_1470,
     csa_tree_add_69_2_groupi_n_1471, csa_tree_add_69_2_groupi_n_1472,
     csa_tree_add_69_2_groupi_n_1473, csa_tree_add_69_2_groupi_n_1474,
     csa_tree_add_69_2_groupi_n_1475, csa_tree_add_69_2_groupi_n_1476,
     csa_tree_add_69_2_groupi_n_1477, csa_tree_add_69_2_groupi_n_1478,
     csa_tree_add_69_2_groupi_n_1479, csa_tree_add_69_2_groupi_n_1481,
     csa_tree_add_69_2_groupi_n_1482, csa_tree_add_69_2_groupi_n_1483,
     csa_tree_add_69_2_groupi_n_1484, csa_tree_add_69_2_groupi_n_1485,
     csa_tree_add_69_2_groupi_n_1486, csa_tree_add_69_2_groupi_n_1487,
     csa_tree_add_69_2_groupi_n_1488, csa_tree_add_69_2_groupi_n_1489,
     csa_tree_add_69_2_groupi_n_1490, csa_tree_add_69_2_groupi_n_1491,
     csa_tree_add_69_2_groupi_n_1492, csa_tree_add_69_2_groupi_n_1493,
     csa_tree_add_69_2_groupi_n_1494, csa_tree_add_69_2_groupi_n_1495,
     csa_tree_add_69_2_groupi_n_1496, csa_tree_add_69_2_groupi_n_1497,
     csa_tree_add_69_2_groupi_n_1498, csa_tree_add_69_2_groupi_n_1499,
     csa_tree_add_69_2_groupi_n_1500, csa_tree_add_69_2_groupi_n_1501,
     csa_tree_add_69_2_groupi_n_1502, csa_tree_add_69_2_groupi_n_1503,
     csa_tree_add_69_2_groupi_n_1504, csa_tree_add_69_2_groupi_n_1505,
     csa_tree_add_69_2_groupi_n_1506, csa_tree_add_69_2_groupi_n_1507,
     csa_tree_add_69_2_groupi_n_1508, csa_tree_add_69_2_groupi_n_1509,
     csa_tree_add_69_2_groupi_n_1510, csa_tree_add_69_2_groupi_n_1511,
     csa_tree_add_69_2_groupi_n_1512, csa_tree_add_69_2_groupi_n_1513,
     csa_tree_add_69_2_groupi_n_1514, csa_tree_add_69_2_groupi_n_1515,
     csa_tree_add_69_2_groupi_n_1516, csa_tree_add_69_2_groupi_n_1517,
     csa_tree_add_69_2_groupi_n_1518, csa_tree_add_69_2_groupi_n_1519,
     csa_tree_add_69_2_groupi_n_1520, csa_tree_add_69_2_groupi_n_1521,
     csa_tree_add_69_2_groupi_n_1522, csa_tree_add_69_2_groupi_n_1523,
     csa_tree_add_69_2_groupi_n_1524, csa_tree_add_69_2_groupi_n_1525,
     csa_tree_add_69_2_groupi_n_1526, csa_tree_add_69_2_groupi_n_1527,
     csa_tree_add_69_2_groupi_n_1528, csa_tree_add_69_2_groupi_n_1529,
     csa_tree_add_69_2_groupi_n_1530, csa_tree_add_69_2_groupi_n_1531,
     csa_tree_add_69_2_groupi_n_1532, csa_tree_add_69_2_groupi_n_1533,
     csa_tree_add_69_2_groupi_n_1534, csa_tree_add_69_2_groupi_n_1535,
     csa_tree_add_69_2_groupi_n_1536, csa_tree_add_69_2_groupi_n_1537,
     csa_tree_add_69_2_groupi_n_1538, csa_tree_add_69_2_groupi_n_1539,
     csa_tree_add_69_2_groupi_n_1540, csa_tree_add_69_2_groupi_n_1541,
     csa_tree_add_69_2_groupi_n_1542, csa_tree_add_69_2_groupi_n_1543,
     csa_tree_add_69_2_groupi_n_1548, csa_tree_add_69_2_groupi_n_1555,
     csa_tree_add_69_2_groupi_n_1556, csa_tree_add_69_2_groupi_n_1557,
     csa_tree_add_69_2_groupi_n_1560, csa_tree_add_69_2_groupi_n_1561,
     csa_tree_add_69_2_groupi_n_1562, csa_tree_add_69_2_groupi_n_1563,
     csa_tree_add_69_2_groupi_n_1564, csa_tree_add_69_2_groupi_n_1565,
     csa_tree_add_69_2_groupi_n_1567, csa_tree_add_69_2_groupi_n_1581,
     csa_tree_add_69_2_groupi_n_1582, csa_tree_add_69_2_groupi_n_1583,
     mul_72_11_n_0, mul_72_11_n_1, mul_72_11_n_2, mul_72_11_n_3, mul_72_11_n_10,
     mul_72_11_n_11, mul_72_11_n_12, mul_72_11_n_13, mul_72_11_n_14,
     mul_72_11_n_15, mul_72_11_n_24, mul_72_11_n_28, mul_72_11_n_37,
     mul_72_11_n_38, mul_72_11_n_39, mul_72_11_n_44, mul_72_11_n_45,
     mul_72_11_n_46, mul_72_11_n_47, mul_72_11_n_49, mul_72_11_n_55,
     mul_72_11_n_59, mul_72_11_n_60, mul_72_11_n_61, mul_72_11_n_62,
     mul_72_11_n_63, mul_72_11_n_66, mul_72_11_n_67, mul_72_11_n_68,
     mul_72_11_n_69, mul_72_11_n_70, mul_72_11_n_71, mul_72_11_n_72,
     mul_72_11_n_73, mul_72_11_n_74, mul_72_11_n_75, mul_72_11_n_76,
     mul_72_11_n_77, mul_72_11_n_79, mul_72_11_n_80, mul_72_11_n_81,
     mul_72_11_n_82, mul_72_11_n_83, mul_72_11_n_84, mul_72_11_n_85,
     mul_72_11_n_86, mul_72_11_n_87, mul_72_11_n_88, mul_72_11_n_89,
     mul_72_11_n_90, mul_72_11_n_91, mul_72_11_n_92, mul_72_11_n_93,
     mul_72_11_n_94, mul_72_11_n_95, mul_72_11_n_96, mul_72_11_n_97,
     mul_72_11_n_98, mul_72_11_n_99, mul_72_11_n_100, mul_72_11_n_101,
     mul_72_11_n_102, mul_72_11_n_103, mul_72_11_n_104, mul_72_11_n_105,
     mul_72_11_n_106, mul_72_11_n_107, mul_72_11_n_108, mul_72_11_n_109,
     mul_72_11_n_110, mul_72_11_n_111, mul_72_11_n_112, mul_72_11_n_113,
     mul_72_11_n_114, mul_72_11_n_115, mul_72_11_n_116, mul_72_11_n_117,
     mul_72_11_n_118, mul_72_11_n_119, mul_72_11_n_120, mul_72_11_n_121,
     mul_72_11_n_122, mul_72_11_n_123, mul_72_11_n_124, mul_72_11_n_125,
     mul_72_11_n_126, mul_72_11_n_127, mul_72_11_n_128, mul_72_11_n_129,
     mul_72_11_n_130, mul_72_11_n_131, mul_72_11_n_132, mul_72_11_n_133,
     mul_72_11_n_134, mul_72_11_n_135, mul_72_11_n_136, mul_72_11_n_137,
     mul_72_11_n_138, mul_72_11_n_139, mul_72_11_n_140, mul_72_11_n_141,
     mul_72_11_n_142, mul_72_11_n_143, mul_72_11_n_144, mul_72_11_n_145,
     mul_72_11_n_146, mul_72_11_n_147, mul_72_11_n_148, mul_72_11_n_149,
     mul_72_11_n_150, mul_72_11_n_151, mul_72_11_n_152, mul_72_11_n_153,
     mul_72_11_n_154, mul_72_11_n_155, mul_72_11_n_156, mul_72_11_n_157,
     mul_72_11_n_158, mul_72_11_n_159, mul_72_11_n_160, mul_72_11_n_161,
     mul_72_11_n_162, mul_72_11_n_163, mul_72_11_n_164, mul_72_11_n_165,
     mul_72_11_n_166, mul_72_11_n_167, mul_72_11_n_168, mul_72_11_n_169,
     mul_72_11_n_170, mul_72_11_n_171, mul_72_11_n_172, mul_72_11_n_173,
     mul_72_11_n_174, mul_72_11_n_175, mul_72_11_n_176, mul_72_11_n_177,
     mul_72_11_n_178, mul_72_11_n_179, mul_72_11_n_180, mul_72_11_n_181,
     mul_72_11_n_182, mul_72_11_n_183, mul_72_11_n_184, mul_72_11_n_185,
     mul_72_11_n_186, mul_72_11_n_187, mul_72_11_n_188, mul_72_11_n_189,
     mul_72_11_n_190, mul_72_11_n_191, mul_72_11_n_192, mul_72_11_n_193,
     mul_72_11_n_194, mul_72_11_n_195, mul_72_11_n_196, mul_72_11_n_197,
     mul_72_11_n_198, mul_72_11_n_199, mul_72_11_n_200, mul_72_11_n_201,
     mul_72_11_n_202, mul_72_11_n_203, mul_72_11_n_204, mul_72_11_n_205,
     mul_72_11_n_206, mul_72_11_n_207, mul_72_11_n_208, mul_72_11_n_209,
     mul_72_11_n_210, mul_72_11_n_211, mul_72_11_n_212, mul_72_11_n_213,
     mul_72_11_n_214, mul_72_11_n_215, mul_72_11_n_216, mul_72_11_n_217,
     mul_72_11_n_218, mul_72_11_n_219, mul_72_11_n_221, mul_72_11_n_222,
     mul_72_11_n_223, mul_72_11_n_224, mul_72_11_n_225, mul_72_11_n_226,
     mul_72_11_n_227, mul_72_11_n_228, mul_72_11_n_229, mul_72_11_n_230,
     mul_72_11_n_231, mul_72_11_n_232, mul_72_11_n_233, mul_72_11_n_234,
     mul_72_11_n_235, mul_72_11_n_236, mul_72_11_n_237, mul_72_11_n_238,
     mul_72_11_n_239, mul_72_11_n_240, mul_72_11_n_241, mul_72_11_n_242,
     mul_72_11_n_243, mul_72_11_n_244, mul_72_11_n_245, mul_72_11_n_246,
     mul_72_11_n_247, mul_72_11_n_248, mul_72_11_n_249, mul_72_11_n_250,
     mul_72_11_n_251, mul_72_11_n_252, mul_72_11_n_253, mul_72_11_n_254,
     mul_72_11_n_255, mul_72_11_n_256, mul_72_11_n_257, mul_72_11_n_258,
     mul_72_11_n_259, mul_72_11_n_260, mul_72_11_n_261, mul_72_11_n_262,
     mul_72_11_n_263, mul_72_11_n_264, mul_72_11_n_265, mul_72_11_n_266,
     mul_72_11_n_267, mul_72_11_n_268, mul_72_11_n_269, mul_72_11_n_270,
     mul_72_11_n_271, mul_72_11_n_272, mul_72_11_n_273, mul_72_11_n_274,
     mul_72_11_n_275, mul_72_11_n_276, mul_72_11_n_277, mul_72_11_n_278,
     mul_72_11_n_279, mul_72_11_n_280, mul_72_11_n_281, mul_72_11_n_282,
     mul_72_11_n_283, mul_72_11_n_284, mul_72_11_n_285, mul_72_11_n_286,
     mul_72_11_n_287, mul_72_11_n_288, mul_72_11_n_289, mul_72_11_n_290,
     mul_72_11_n_291, mul_72_11_n_292, mul_72_11_n_293, mul_72_11_n_294,
     mul_72_11_n_295, mul_72_11_n_296, mul_72_11_n_297, mul_72_11_n_298,
     mul_72_11_n_299, mul_72_11_n_300, mul_72_11_n_301, mul_72_11_n_302,
     mul_72_11_n_303, mul_72_11_n_304, mul_72_11_n_305, mul_72_11_n_306,
     mul_72_11_n_307, mul_72_11_n_308, mul_72_11_n_309, mul_72_11_n_310,
     mul_72_11_n_311, mul_72_11_n_312, mul_72_11_n_313, mul_72_11_n_314,
     mul_72_11_n_315, mul_72_11_n_316, mul_72_11_n_317, mul_72_11_n_318,
     mul_72_11_n_319, mul_72_11_n_320, mul_72_11_n_321, mul_72_11_n_322,
     mul_72_11_n_323, mul_72_11_n_324, mul_72_11_n_325, mul_72_11_n_326,
     mul_72_11_n_327, mul_72_11_n_328, mul_72_11_n_329, mul_72_11_n_330,
     mul_72_11_n_331, mul_72_11_n_332, mul_72_11_n_333, mul_72_11_n_334,
     mul_72_11_n_335, mul_72_11_n_336, mul_72_11_n_337, mul_72_11_n_338,
     mul_72_11_n_339, mul_72_11_n_340, mul_72_11_n_341, mul_72_11_n_342,
     mul_72_11_n_343, mul_72_11_n_344, mul_72_11_n_345, mul_72_11_n_346,
     mul_72_11_n_347, mul_72_11_n_348, mul_72_11_n_349, mul_72_11_n_350,
     mul_72_11_n_351, mul_72_11_n_352, mul_72_11_n_353, mul_72_11_n_354,
     mul_72_11_n_355, mul_72_11_n_356, mul_72_11_n_357, mul_72_11_n_358,
     mul_72_11_n_359, mul_72_11_n_360, mul_72_11_n_361, mul_72_11_n_362,
     mul_72_11_n_363, mul_72_11_n_364, mul_72_11_n_365, mul_72_11_n_366,
     mul_72_11_n_367, mul_72_11_n_368, mul_72_11_n_369, mul_72_11_n_370,
     mul_72_11_n_371, mul_72_11_n_372, mul_72_11_n_373, mul_72_11_n_374,
     mul_72_11_n_375, mul_72_11_n_376, mul_72_11_n_377, mul_72_11_n_378,
     mul_72_11_n_379, mul_72_11_n_380, mul_72_11_n_381, mul_72_11_n_382,
     mul_72_11_n_383, mul_72_11_n_384, mul_72_11_n_385, mul_72_11_n_386,
     mul_72_11_n_387, mul_72_11_n_388, mul_72_11_n_389, mul_72_11_n_390,
     mul_72_11_n_391, mul_72_11_n_392, mul_72_11_n_393, mul_72_11_n_394,
     mul_72_11_n_395, mul_72_11_n_396, mul_72_11_n_397, mul_72_11_n_398,
     mul_72_11_n_399, mul_72_11_n_400, mul_72_11_n_401, mul_72_11_n_402,
     mul_72_11_n_403, mul_72_11_n_404, mul_72_11_n_405, mul_72_11_n_406,
     mul_72_11_n_407, mul_72_11_n_408, mul_72_11_n_409, mul_72_11_n_410,
     mul_72_11_n_411, mul_72_11_n_412, mul_72_11_n_413, mul_72_11_n_414,
     mul_72_11_n_415, mul_72_11_n_416, mul_72_11_n_417, mul_72_11_n_418,
     mul_72_11_n_419, mul_72_11_n_420, mul_72_11_n_421, mul_72_11_n_422,
     mul_72_11_n_423, mul_72_11_n_424, mul_72_11_n_425, mul_72_11_n_426,
     mul_72_11_n_427, mul_72_11_n_428, mul_72_11_n_429, mul_72_11_n_430,
     mul_72_11_n_431, mul_72_11_n_432, mul_72_11_n_433, mul_72_11_n_434,
     mul_72_11_n_435, mul_72_11_n_436, mul_72_11_n_437, mul_72_11_n_438,
     mul_72_11_n_439, mul_72_11_n_440, mul_72_11_n_441, mul_72_11_n_442,
     mul_72_11_n_443, mul_72_11_n_444, mul_72_11_n_445, mul_72_11_n_446,
     mul_72_11_n_447, mul_72_11_n_448, mul_72_11_n_449, mul_72_11_n_450,
     mul_72_11_n_451, mul_72_11_n_452, mul_72_11_n_453, mul_72_11_n_454,
     mul_72_11_n_455, mul_72_11_n_456, mul_72_11_n_457, mul_72_11_n_458,
     mul_72_11_n_459, mul_72_11_n_460, mul_72_11_n_461, mul_72_11_n_462,
     mul_72_11_n_463, mul_72_11_n_464, mul_72_11_n_465, mul_72_11_n_466,
     mul_72_11_n_467, mul_72_11_n_468, mul_72_11_n_469, mul_72_11_n_470,
     mul_72_11_n_471, mul_72_11_n_472, mul_72_11_n_473, mul_72_11_n_474,
     mul_72_11_n_475, mul_72_11_n_476, mul_72_11_n_477, mul_72_11_n_478,
     mul_72_11_n_479, mul_72_11_n_480, mul_72_11_n_481, mul_72_11_n_482,
     mul_72_11_n_483, mul_72_11_n_484, mul_72_11_n_485, mul_72_11_n_486,
     mul_72_11_n_487, mul_72_11_n_488, mul_72_11_n_489, mul_72_11_n_490,
     mul_72_11_n_491, mul_72_11_n_492, mul_72_11_n_493, mul_72_11_n_494,
     mul_72_11_n_495, mul_72_11_n_496, mul_72_11_n_497, mul_72_11_n_498,
     mul_72_11_n_499, mul_72_11_n_500, mul_72_11_n_501, mul_72_11_n_502,
     mul_72_11_n_503, mul_72_11_n_504, mul_72_11_n_505, mul_72_11_n_506,
     mul_72_11_n_507, mul_72_11_n_508, mul_72_11_n_509, mul_72_11_n_510,
     mul_72_11_n_511, mul_72_11_n_512, mul_72_11_n_513, mul_72_11_n_514,
     mul_72_11_n_515, mul_72_11_n_516, mul_72_11_n_517, mul_72_11_n_518,
     mul_72_11_n_519, mul_72_11_n_520, mul_72_11_n_521, mul_72_11_n_522,
     mul_72_11_n_523, mul_72_11_n_524, mul_72_11_n_525, mul_72_11_n_526,
     mul_72_11_n_527, mul_72_11_n_528, mul_72_11_n_529, mul_72_11_n_530,
     mul_72_11_n_531, mul_72_11_n_532, mul_72_11_n_533, mul_72_11_n_534,
     mul_72_11_n_535, mul_72_11_n_536, mul_72_11_n_537, mul_72_11_n_538,
     mul_72_11_n_539, mul_72_11_n_540, mul_72_11_n_541, mul_72_11_n_542,
     mul_72_11_n_543, mul_72_11_n_544, mul_72_11_n_545, mul_72_11_n_546,
     mul_72_11_n_547, mul_72_11_n_548, mul_72_11_n_549, mul_72_11_n_550,
     mul_72_11_n_551, mul_72_11_n_552, mul_72_11_n_553, mul_72_11_n_554,
     mul_72_11_n_555, mul_72_11_n_556, mul_72_11_n_557, mul_72_11_n_558,
     mul_72_11_n_559, mul_72_11_n_560, mul_72_11_n_561, mul_72_11_n_562,
     mul_72_11_n_563, mul_72_11_n_564, mul_72_11_n_565, mul_72_11_n_566,
     mul_72_11_n_567, mul_72_11_n_568, mul_72_11_n_569, mul_72_11_n_570,
     mul_72_11_n_571, mul_72_11_n_572, mul_72_11_n_573, mul_72_11_n_574,
     mul_72_11_n_575, mul_72_11_n_576, mul_72_11_n_577, mul_72_11_n_578,
     mul_72_11_n_579, mul_72_11_n_580, mul_72_11_n_581, mul_72_11_n_582,
     mul_72_11_n_583, mul_72_11_n_584, mul_72_11_n_585, mul_72_11_n_586,
     mul_72_11_n_587, mul_72_11_n_588, mul_72_11_n_589, mul_72_11_n_590,
     mul_72_11_n_591, mul_72_11_n_592, mul_72_11_n_593, mul_72_11_n_594,
     mul_72_11_n_595, mul_72_11_n_596, mul_72_11_n_597, mul_72_11_n_598,
     mul_72_11_n_599, mul_72_11_n_600, mul_72_11_n_601, mul_72_11_n_602,
     mul_72_11_n_603, mul_72_11_n_604, mul_72_11_n_605, mul_72_11_n_606,
     mul_72_11_n_607, mul_72_11_n_608, mul_72_11_n_609, mul_72_11_n_610,
     mul_72_11_n_611, mul_72_11_n_612, mul_72_11_n_613, mul_72_11_n_614,
     mul_72_11_n_615, mul_72_11_n_616, mul_72_11_n_617, mul_72_11_n_618,
     mul_72_11_n_619, mul_72_11_n_620, mul_72_11_n_621, mul_72_11_n_622,
     mul_72_11_n_623, mul_72_11_n_624, mul_72_11_n_625, mul_72_11_n_626,
     mul_72_11_n_627, mul_72_11_n_628, mul_72_11_n_629, mul_72_11_n_630,
     mul_72_11_n_631, mul_72_11_n_632, mul_72_11_n_633, mul_72_11_n_634,
     mul_72_11_n_635, mul_72_11_n_636, mul_72_11_n_637, mul_72_11_n_638,
     mul_72_11_n_639, mul_72_11_n_640, mul_72_11_n_641, mul_72_11_n_642,
     mul_72_11_n_643, mul_72_11_n_644, mul_72_11_n_645, mul_72_11_n_646,
     mul_72_11_n_647, mul_72_11_n_648, mul_72_11_n_649, mul_72_11_n_650,
     mul_72_11_n_651, mul_72_11_n_652, mul_72_11_n_653, mul_72_11_n_654,
     mul_72_11_n_655, mul_72_11_n_656, mul_72_11_n_657, mul_72_11_n_658,
     mul_72_11_n_659, mul_72_11_n_660, mul_72_11_n_661, mul_72_11_n_662,
     mul_72_11_n_663, mul_72_11_n_664, mul_72_11_n_665, mul_72_11_n_666,
     mul_72_11_n_667, mul_72_11_n_668, mul_72_11_n_669, mul_72_11_n_670,
     mul_72_11_n_671, mul_72_11_n_672, mul_72_11_n_673, mul_72_11_n_674,
     mul_72_11_n_675, mul_72_11_n_676, mul_72_11_n_677, mul_72_11_n_678,
     mul_72_11_n_679, mul_72_11_n_680, mul_72_11_n_681, mul_72_11_n_682,
     mul_72_11_n_683, mul_72_11_n_684, mul_72_11_n_685, mul_72_11_n_686,
     mul_72_11_n_687, mul_72_11_n_688, mul_72_11_n_689, mul_72_11_n_690,
     mul_72_11_n_692, mul_72_11_n_693, mul_72_11_n_694, mul_72_11_n_695,
     mul_72_11_n_696, mul_72_11_n_697, mul_72_11_n_698, mul_72_11_n_699,
     mul_72_11_n_700, mul_72_11_n_701, mul_72_11_n_702, mul_72_11_n_703,
     mul_72_11_n_704, mul_72_11_n_705, mul_72_11_n_706, mul_72_11_n_707,
     mul_72_11_n_708, mul_72_11_n_709, mul_72_11_n_710, mul_72_11_n_711,
     mul_72_11_n_712, mul_72_11_n_713, mul_72_11_n_714, mul_72_11_n_715,
     mul_72_11_n_716, mul_72_11_n_717, mul_72_11_n_718, mul_72_11_n_719,
     mul_72_11_n_720, mul_72_11_n_721, mul_72_11_n_722, mul_72_11_n_723,
     mul_72_11_n_724, mul_72_11_n_725, mul_72_11_n_726, mul_72_11_n_727,
     mul_72_11_n_728, mul_72_11_n_729, mul_72_11_n_730, mul_72_11_n_731,
     mul_72_11_n_732, mul_72_11_n_733, mul_72_11_n_734, mul_72_11_n_735,
     mul_72_11_n_736, mul_72_11_n_737, mul_72_11_n_738, mul_72_11_n_739,
     mul_72_11_n_740, mul_72_11_n_741, mul_72_11_n_742, mul_72_11_n_743,
     mul_72_11_n_744, mul_72_11_n_745, mul_72_11_n_746, mul_72_11_n_748,
     mul_72_11_n_749, mul_72_11_n_750, mul_72_11_n_751, mul_72_11_n_752,
     mul_72_11_n_753, mul_72_11_n_754, mul_72_11_n_755, mul_72_11_n_756,
     mul_72_11_n_757, mul_72_11_n_758, mul_72_11_n_759, mul_72_11_n_760,
     mul_72_11_n_761, mul_72_11_n_762, mul_72_11_n_763, mul_72_11_n_764,
     mul_72_11_n_765, mul_72_11_n_766, mul_72_11_n_767, mul_72_11_n_768,
     mul_72_11_n_769, mul_72_11_n_770, mul_72_11_n_771, mul_72_11_n_772,
     mul_72_11_n_773, mul_72_11_n_774, mul_72_11_n_775, mul_72_11_n_776,
     mul_72_11_n_777, mul_72_11_n_778, mul_72_11_n_779, mul_72_11_n_780,
     mul_72_11_n_781, mul_72_11_n_782, mul_72_11_n_783, mul_72_11_n_784,
     mul_72_11_n_785, mul_72_11_n_786, mul_72_11_n_787, mul_72_11_n_788,
     mul_72_11_n_789, mul_72_11_n_790, mul_72_11_n_791, mul_72_11_n_792,
     mul_72_11_n_793, mul_72_11_n_794, mul_72_11_n_795, mul_72_11_n_796,
     mul_72_11_n_797, mul_72_11_n_798, mul_72_11_n_799, mul_72_11_n_800,
     mul_72_11_n_801, mul_72_11_n_802, mul_72_11_n_803, mul_72_11_n_804,
     mul_72_11_n_805, mul_72_11_n_806, mul_72_11_n_807, mul_72_11_n_808,
     mul_72_11_n_810, mul_72_11_n_811, mul_72_11_n_812, mul_72_11_n_813,
     mul_72_11_n_814, mul_72_11_n_815, mul_72_11_n_816, mul_72_11_n_817,
     mul_72_11_n_818, mul_72_11_n_819, mul_72_11_n_820, mul_72_11_n_821,
     mul_72_11_n_822, mul_72_11_n_823, mul_72_11_n_824, mul_72_11_n_825,
     mul_72_11_n_826, mul_72_11_n_827, mul_72_11_n_828, mul_72_11_n_829,
     mul_72_11_n_830, mul_72_11_n_831, mul_72_11_n_832, mul_72_11_n_833,
     mul_72_11_n_834, mul_72_11_n_835, mul_72_11_n_836, mul_72_11_n_837,
     mul_72_11_n_838, mul_72_11_n_839, mul_72_11_n_840, mul_72_11_n_841,
     mul_72_11_n_842, mul_72_11_n_843, mul_72_11_n_844, mul_72_11_n_845,
     mul_72_11_n_846, mul_72_11_n_847, mul_72_11_n_848, mul_72_11_n_849,
     mul_72_11_n_850, mul_72_11_n_851, mul_72_11_n_852, mul_72_11_n_853,
     mul_72_11_n_854, mul_72_11_n_855, mul_72_11_n_857, mul_72_11_n_858,
     mul_72_11_n_859, mul_72_11_n_860, mul_72_11_n_861, mul_72_11_n_862,
     mul_72_11_n_863, mul_72_11_n_864, mul_72_11_n_865, mul_72_11_n_866,
     mul_72_11_n_867, mul_72_11_n_868, mul_72_11_n_869, mul_72_11_n_870,
     mul_72_11_n_871, mul_72_11_n_872, mul_72_11_n_873, mul_72_11_n_874,
     mul_72_11_n_875, mul_72_11_n_876, mul_72_11_n_877, mul_72_11_n_878,
     mul_72_11_n_879, mul_72_11_n_880, mul_72_11_n_881, mul_72_11_n_882,
     mul_72_11_n_883, mul_72_11_n_884, mul_72_11_n_885, mul_72_11_n_886,
     mul_72_11_n_887, mul_72_11_n_888, mul_72_11_n_889, mul_72_11_n_890,
     mul_72_11_n_891, mul_72_11_n_892, mul_72_11_n_893, mul_72_11_n_894,
     mul_72_11_n_895, mul_72_11_n_896, mul_72_11_n_897, mul_72_11_n_898,
     mul_72_11_n_899, mul_72_11_n_900, mul_72_11_n_901, mul_72_11_n_903,
     mul_72_11_n_904, mul_72_11_n_905, mul_72_11_n_906, mul_72_11_n_907,
     mul_72_11_n_908, mul_72_11_n_909, mul_72_11_n_910, mul_72_11_n_911,
     mul_72_11_n_912, mul_72_11_n_913, mul_72_11_n_914, mul_72_11_n_915,
     mul_72_11_n_916, mul_72_11_n_917, mul_72_11_n_918, mul_72_11_n_919,
     mul_72_11_n_920, mul_72_11_n_921, mul_72_11_n_922, mul_72_11_n_923,
     mul_72_11_n_924, mul_72_11_n_925, mul_72_11_n_926, mul_72_11_n_927,
     mul_72_11_n_928, mul_72_11_n_929, mul_72_11_n_930, mul_72_11_n_931,
     mul_72_11_n_932, mul_72_11_n_933, mul_72_11_n_934, mul_72_11_n_935,
     mul_72_11_n_936, mul_72_11_n_937, mul_72_11_n_938, mul_72_11_n_939,
     mul_72_11_n_940, mul_72_11_n_941, mul_72_11_n_943, mul_72_11_n_944,
     mul_72_11_n_945, mul_72_11_n_946, mul_72_11_n_947, mul_72_11_n_948,
     mul_72_11_n_949, mul_72_11_n_950, mul_72_11_n_951, mul_72_11_n_952,
     mul_72_11_n_953, mul_72_11_n_954, mul_72_11_n_955, mul_72_11_n_956,
     mul_72_11_n_957, mul_72_11_n_958, mul_72_11_n_959, mul_72_11_n_960,
     mul_72_11_n_961, mul_72_11_n_962, mul_72_11_n_963, mul_72_11_n_964,
     mul_72_11_n_965, mul_72_11_n_966, mul_72_11_n_967, mul_72_11_n_968,
     mul_72_11_n_969, mul_72_11_n_970, mul_72_11_n_971, mul_72_11_n_972,
     mul_72_11_n_973, mul_72_11_n_974, mul_72_11_n_975, mul_72_11_n_976,
     mul_72_11_n_977, mul_72_11_n_978, mul_72_11_n_979, mul_72_11_n_980,
     mul_72_11_n_981, mul_72_11_n_982, mul_72_11_n_983, mul_72_11_n_984,
     mul_72_11_n_985, mul_72_11_n_986, mul_72_11_n_988, mul_72_11_n_989,
     mul_72_11_n_990, mul_72_11_n_991, mul_72_11_n_992, mul_72_11_n_993,
     mul_72_11_n_994, mul_72_11_n_995, mul_72_11_n_996, mul_72_11_n_997,
     mul_72_11_n_998, mul_72_11_n_999, mul_72_11_n_1000, mul_72_11_n_1001,
     mul_72_11_n_1002, mul_72_11_n_1003, mul_72_11_n_1004, mul_72_11_n_1005,
     mul_72_11_n_1006, mul_72_11_n_1007, mul_72_11_n_1008, mul_72_11_n_1009,
     mul_72_11_n_1010, mul_72_11_n_1011, mul_72_11_n_1012, mul_72_11_n_1013,
     mul_72_11_n_1014, mul_72_11_n_1015, mul_72_11_n_1016, mul_72_11_n_1017,
     mul_72_11_n_1018, mul_72_11_n_1019, mul_72_11_n_1020, mul_72_11_n_1021,
     mul_72_11_n_1022, mul_72_11_n_1023, mul_72_11_n_1024, mul_72_11_n_1025,
     mul_72_11_n_1026, mul_72_11_n_1027, mul_72_11_n_1028, mul_72_11_n_1029,
     mul_72_11_n_1030, mul_72_11_n_1031, mul_72_11_n_1032, mul_72_11_n_1033,
     mul_72_11_n_1034, mul_72_11_n_1035, mul_72_11_n_1036, mul_72_11_n_1037,
     mul_72_11_n_1038, mul_72_11_n_1039, mul_72_11_n_1040, mul_72_11_n_1041,
     mul_72_11_n_1042, mul_72_11_n_1043, mul_72_11_n_1045, mul_72_11_n_1046,
     mul_72_11_n_1047, mul_72_11_n_1048, mul_72_11_n_1049, mul_72_11_n_1050,
     mul_72_11_n_1051, mul_72_11_n_1052, mul_72_11_n_1053, mul_72_11_n_1054,
     mul_72_11_n_1055, mul_72_11_n_1056, mul_72_11_n_1057, mul_72_11_n_1058,
     mul_72_11_n_1059, mul_72_11_n_1060, mul_72_11_n_1061, mul_72_11_n_1062,
     mul_72_11_n_1063, mul_72_11_n_1064, mul_72_11_n_1065, mul_72_11_n_1066,
     mul_72_11_n_1067, mul_72_11_n_1068, mul_72_11_n_1069, mul_72_11_n_1070,
     mul_72_11_n_1071, mul_72_11_n_1072, mul_72_11_n_1073, mul_72_11_n_1074,
     mul_72_11_n_1075, mul_72_11_n_1076, mul_72_11_n_1077, mul_72_11_n_1078,
     mul_72_11_n_1079, mul_72_11_n_1080, mul_72_11_n_1081, mul_72_11_n_1082,
     mul_72_11_n_1083, mul_72_11_n_1084, mul_72_11_n_1085, mul_72_11_n_1088,
     mul_72_11_n_1089, mul_72_11_n_1090, mul_72_11_n_1091, mul_72_11_n_1092,
     mul_72_11_n_1093, mul_72_11_n_1094, mul_72_11_n_1095, mul_72_11_n_1096,
     mul_72_11_n_1097, mul_72_11_n_1098, mul_72_11_n_1099, mul_72_11_n_1100,
     mul_72_11_n_1101, mul_72_11_n_1102, mul_72_11_n_1103, mul_72_11_n_1104,
     mul_72_11_n_1105, mul_72_11_n_1106, mul_72_11_n_1107, mul_72_11_n_1108,
     mul_72_11_n_1109, mul_72_11_n_1110, mul_72_11_n_1111, mul_72_11_n_1112,
     mul_72_11_n_1113, mul_72_11_n_1114, mul_72_11_n_1115, mul_72_11_n_1116,
     mul_72_11_n_1117, mul_72_11_n_1119, mul_72_11_n_1120, mul_72_11_n_1121,
     mul_72_11_n_1122, mul_72_11_n_1123, mul_72_11_n_1124, mul_72_11_n_1125,
     mul_72_11_n_1126, mul_72_11_n_1127, mul_72_11_n_1128, mul_72_11_n_1129,
     mul_72_11_n_1130, mul_72_11_n_1131, mul_72_11_n_1132, mul_72_11_n_1133,
     mul_72_11_n_1134, mul_72_11_n_1135, mul_72_11_n_1136, mul_72_11_n_1137,
     mul_72_11_n_1138, mul_72_11_n_1139, mul_72_11_n_1140, mul_72_11_n_1141,
     mul_72_11_n_1142, mul_72_11_n_1143, mul_72_11_n_1144, mul_72_11_n_1145,
     mul_72_11_n_1146, mul_72_11_n_1147, mul_72_11_n_1148, mul_72_11_n_1149,
     mul_72_11_n_1150, mul_72_11_n_1151, mul_72_11_n_1152, mul_72_11_n_1153,
     mul_72_11_n_1154, mul_72_11_n_1155, mul_72_11_n_1156, mul_72_11_n_1157,
     mul_72_11_n_1158, mul_72_11_n_1159, mul_72_11_n_1161, mul_72_11_n_1162,
     mul_72_11_n_1163, mul_72_11_n_1164, mul_72_11_n_1165, mul_72_11_n_1166,
     mul_72_11_n_1167, mul_72_11_n_1168, mul_72_11_n_1169, mul_72_11_n_1170,
     mul_72_11_n_1171, mul_72_11_n_1172, mul_72_11_n_1173, mul_72_11_n_1174,
     mul_72_11_n_1175, mul_72_11_n_1176, mul_72_11_n_1177, mul_72_11_n_1178,
     mul_72_11_n_1179, mul_72_11_n_1180, mul_72_11_n_1181, mul_72_11_n_1182,
     mul_72_11_n_1183, mul_72_11_n_1184, mul_72_11_n_1185, mul_72_11_n_1186,
     mul_72_11_n_1187, mul_72_11_n_1188, mul_72_11_n_1189, mul_72_11_n_1190,
     mul_72_11_n_1193, mul_72_11_n_1194, mul_72_11_n_1195, mul_72_11_n_1196,
     mul_72_11_n_1197, mul_72_11_n_1198, mul_72_11_n_1199, mul_72_11_n_1200,
     mul_72_11_n_1201, mul_72_11_n_1202, mul_72_11_n_1203, mul_72_11_n_1204,
     mul_72_11_n_1205, mul_72_11_n_1206, mul_72_11_n_1207, mul_72_11_n_1208,
     mul_72_11_n_1209, mul_72_11_n_1210, mul_72_11_n_1211, mul_72_11_n_1212,
     mul_72_11_n_1213, mul_72_11_n_1215, mul_72_11_n_1216, mul_72_11_n_1217,
     mul_72_11_n_1218, mul_72_11_n_1219, mul_72_11_n_1220, mul_72_11_n_1221,
     mul_72_11_n_1222, mul_72_11_n_1223, mul_72_11_n_1224, mul_72_11_n_1225,
     mul_72_11_n_1226, mul_72_11_n_1227, mul_72_11_n_1228, mul_72_11_n_1229,
     mul_72_11_n_1230, mul_72_11_n_1231, mul_72_11_n_1232, mul_72_11_n_1233,
     mul_72_11_n_1234, mul_72_11_n_1235, mul_72_11_n_1236, mul_72_11_n_1237,
     mul_72_11_n_1238, mul_72_11_n_1239, mul_72_11_n_1240, mul_72_11_n_1241,
     mul_72_11_n_1242, mul_72_11_n_1243, mul_72_11_n_1244, mul_72_11_n_1245,
     mul_72_11_n_1246, mul_72_11_n_1247, mul_72_11_n_1248, mul_72_11_n_1249,
     mul_72_11_n_1250, mul_72_11_n_1251, mul_72_11_n_1252, mul_72_11_n_1253,
     mul_72_11_n_1254, mul_72_11_n_1255, mul_72_11_n_1256, mul_72_11_n_1257,
     mul_72_11_n_1258, mul_72_11_n_1259, mul_72_11_n_1260, mul_72_11_n_1261,
     mul_72_11_n_1262, mul_72_11_n_1263, mul_72_11_n_1264, mul_72_11_n_1265,
     mul_72_11_n_1266, mul_72_11_n_1267, mul_72_11_n_1268, mul_72_11_n_1269,
     mul_72_11_n_1270, mul_72_11_n_1271, mul_72_11_n_1272, mul_72_11_n_1275,
     mul_72_11_n_1276, mul_72_11_n_1277, mul_72_11_n_1278, mul_72_11_n_1279,
     mul_72_11_n_1280, mul_72_11_n_1281, mul_72_11_n_1282, mul_72_11_n_1283,
     mul_72_11_n_1284, mul_72_11_n_1286, mul_72_11_n_1287, mul_72_11_n_1288,
     mul_72_11_n_1289, mul_72_11_n_1290, mul_72_11_n_1291, mul_72_11_n_1293,
     mul_72_11_n_1296, mul_72_11_n_1297, mul_72_11_n_1298, mul_72_11_n_1301,
     mul_72_11_n_1302, mul_72_11_n_1303, mul_72_11_n_1306, mul_72_11_n_1307,
     mul_72_11_n_1310, mul_72_11_n_1311, mul_72_11_n_1313, mul_72_11_n_1314, n_0,
     n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13, n_14,
     n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25, n_26,
     n_27, n_28, n_29, n_30, n_31, n_32, n_33, n_34, n_35, n_36, n_37, n_38,
     n_39, n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47, n_48, n_49, n_50,
     n_51, n_52, n_53, n_54, n_55, n_56, n_57, n_58, n_59, n_60, n_61, n_62,
     n_63, clk, n_97, n_98, n_99, n_100, n_101, n_102, n_103, n_104, n_105,
     n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113, n_114, n_115, n_116,
     n_117, n_118, n_119, n_120, n_121, n_122, n_123, n_124, n_125, n_126, n_127,
     n_128, n_129, n_130, n_131, n_132, n_133, n_134, n_135, n_136, n_137, n_138,
     n_139, n_140, n_141, n_142, n_143, n_144, n_145, n_146, n_147, n_148, n_149,
     n_150, n_151, n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160,
     n_161, n_162, n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171,
     n_172, n_173, n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182,
     n_183, n_184, n_185, n_186, n_187, n_188, n_189, n_190, n_191, n_192, n_193,
     n_194, n_195, n_196, n_197, n_198, n_199, n_200, n_201, n_202, n_203, n_204,
     n_205, n_206, n_207, n_208, n_209, n_210, n_211, n_212, n_213, n_214, n_215,
     n_216, n_217, n_218, n_219, n_220, n_221, n_222, n_223, n_224, n_225, n_226,
     n_227, n_228, n_229, n_230, n_231, n_232, n_233, n_234, n_235, n_236, n_237,
     n_238, n_239, n_240, n_241, n_242, n_243, n_244, n_245, n_246, n_247, n_248,
     n_249, n_250, n_251, n_252, n_253, n_254, n_255, n_256, n_257, n_258, n_368,
     n_369, n_370, n_371, n_372, n_373, n_374, n_375, n_376, n_377, n_378, n_379,
     n_382, n_388, n_391, n_397, n_398, n_399, n_400, n_401, n_402, n_403, n_404,
     n_405, n_406, n_407, n_408, n_409, n_410, n_411, n_412, n_413, n_414, n_415,
     n_416, n_417, n_418, n_419, n_420, n_421, n_422, n_423, n_424, n_425, n_426,
     n_427, n_428, n_429, n_430, n_431, n_432, n_433, n_434, n_435, n_436, n_437,
     n_438, n_439, n_440, n_441, n_442, n_443, n_444, n_445, n_446, n_447, n_448,
     n_449, n_450, n_451, n_452, n_453, n_454, n_455, n_456, n_457, n_458, n_459,
     n_460, n_461, n_462, n_463, n_464, n_465, n_466, n_467, n_468, n_469, n_470,
     n_471, n_472, n_473, n_474, n_475, n_476, n_477, n_478, n_479, n_480, n_481,
     n_482, n_483, n_484, n_485, n_486, n_487, n_488, n_489, n_490, n_491, n_492,
     n_493, n_494, n_495, n_496, n_497, n_498, n_499, n_500, n_501, n_502, n_503,
     n_504, n_505, n_506, n_507, n_508, n_509, n_510, n_511, n_512, n_513;
 reg retime_s1_1_reg_reg_N30;
 always @(posedge clk)
         retime_s1_1_reg_reg_N30 <= {in3[31]};
 assign n_97 = retime_s1_1_reg_reg_N30;
 reg retime_s1_2_reg_reg_N30;
 always @(posedge clk)
         retime_s1_2_reg_reg_N30 <= n_57;
 assign n_98 = retime_s1_2_reg_reg_N30;
 reg retime_s1_3_reg_reg_N30;
 always @(posedge clk)
         retime_s1_3_reg_reg_N30 <= n_56;
 assign n_99 = retime_s1_3_reg_reg_N30;
 reg retime_s1_4_reg_reg_N30;
 always @(posedge clk)
         retime_s1_4_reg_reg_N30 <= n_38;
 assign n_100 = retime_s1_4_reg_reg_N30;
 reg retime_s1_5_reg_reg_N30;
 always @(posedge clk)
         retime_s1_5_reg_reg_N30 <= n_372;
 assign n_101 = retime_s1_5_reg_reg_N30;
 reg retime_s1_6_reg_reg_N30;
 always @(posedge clk)
         retime_s1_6_reg_reg_N30 <= n_414;
 assign n_102 = retime_s1_6_reg_reg_N30;
 reg retime_s1_7_reg_reg_N30;
 always @(posedge clk)
         retime_s1_7_reg_reg_N30 <= n_419;
 assign n_103 = retime_s1_7_reg_reg_N30;
 reg retime_s1_8_reg_reg_N30;
 always @(posedge clk)
         retime_s1_8_reg_reg_N30 <= n_63;
 assign n_104 = retime_s1_8_reg_reg_N30;
 reg retime_s1_9_reg_reg_N30;
 always @(posedge clk)
         retime_s1_9_reg_reg_N30 <= n_55;
 assign n_105 = retime_s1_9_reg_reg_N30;
 reg retime_s1_10_reg_reg_N30;
 always @(posedge clk)
         retime_s1_10_reg_reg_N30 <= n_43;
 assign n_106 = retime_s1_10_reg_reg_N30;
 reg retime_s1_11_reg_reg_N30;
 always @(posedge clk)
         retime_s1_11_reg_reg_N30 <= n_42;
 assign n_107 = retime_s1_11_reg_reg_N30;
 reg retime_s1_12_reg_reg_N30;
 always @(posedge clk)
         retime_s1_12_reg_reg_N30 <= n_47;
 assign n_108 = retime_s1_12_reg_reg_N30;
 reg retime_s1_13_reg_reg_N30;
 always @(posedge clk)
         retime_s1_13_reg_reg_N30 <= n_46;
 assign n_109 = retime_s1_13_reg_reg_N30;
 reg retime_s1_14_reg_reg_N30;
 always @(posedge clk)
         retime_s1_14_reg_reg_N30 <= n_41;
 assign n_110 = retime_s1_14_reg_reg_N30;
 reg retime_s1_15_reg_reg_N30;
 always @(posedge clk)
         retime_s1_15_reg_reg_N30 <= n_40;
 assign n_111 = retime_s1_15_reg_reg_N30;
 reg retime_s1_16_reg_reg_N30;
 always @(posedge clk)
         retime_s1_16_reg_reg_N30 <= n_51;
 assign n_112 = retime_s1_16_reg_reg_N30;
 reg retime_s1_17_reg_reg_N30;
 always @(posedge clk)
         retime_s1_17_reg_reg_N30 <= n_50;
 assign n_113 = retime_s1_17_reg_reg_N30;
 reg retime_s1_18_reg_reg_N30;
 always @(posedge clk)
         retime_s1_18_reg_reg_N30 <= n_49;
 assign n_114 = retime_s1_18_reg_reg_N30;
 reg retime_s1_19_reg_reg_N30;
 always @(posedge clk)
         retime_s1_19_reg_reg_N30 <= n_48;
 assign n_115 = retime_s1_19_reg_reg_N30;
 reg retime_s1_20_reg_reg_N30;
 always @(posedge clk)
         retime_s1_20_reg_reg_N30 <= n_53;
 assign n_116 = retime_s1_20_reg_reg_N30;
 reg retime_s1_21_reg_reg_N30;
 always @(posedge clk)
         retime_s1_21_reg_reg_N30 <= n_52;
 assign n_117 = retime_s1_21_reg_reg_N30;
 reg retime_s1_22_reg_reg_N30;
 always @(posedge clk)
         retime_s1_22_reg_reg_N30 <= n_37;
 assign n_118 = retime_s1_22_reg_reg_N30;
 reg retime_s1_23_reg_reg_N30;
 always @(posedge clk)
         retime_s1_23_reg_reg_N30 <= n_36;
 assign n_119 = retime_s1_23_reg_reg_N30;
 reg retime_s1_24_reg_reg_N30;
 always @(posedge clk)
         retime_s1_24_reg_reg_N30 <= n_229;
 assign n_120 = retime_s1_24_reg_reg_N30;
 reg retime_s1_25_reg_reg_N30;
 always @(posedge clk)
         retime_s1_25_reg_reg_N30 <= n_45;
 assign n_121 = retime_s1_25_reg_reg_N30;
 reg retime_s1_26_reg_reg_N30;
 always @(posedge clk)
         retime_s1_26_reg_reg_N30 <= n_44;
 assign n_122 = retime_s1_26_reg_reg_N30;
 reg retime_s1_27_reg_reg_N30;
 always @(posedge clk)
         retime_s1_27_reg_reg_N30 <= n_59;
 assign n_123 = retime_s1_27_reg_reg_N30;
 reg retime_s1_28_reg_reg_N30;
 always @(posedge clk)
         retime_s1_28_reg_reg_N30 <= n_58;
 assign n_124 = retime_s1_28_reg_reg_N30;
 reg retime_s1_29_reg_reg_N30;
 always @(posedge clk)
         retime_s1_29_reg_reg_N30 <= n_241;
 assign n_125 = retime_s1_29_reg_reg_N30;
 reg retime_s1_30_reg_reg_N30;
 always @(posedge clk)
         retime_s1_30_reg_reg_N30 <= n_239;
 assign n_126 = retime_s1_30_reg_reg_N30;
 reg retime_s1_31_reg_reg_N30;
 always @(posedge clk)
         retime_s1_31_reg_reg_N30 <= n_222;
 assign n_127 = retime_s1_31_reg_reg_N30;
 reg retime_s1_32_reg_reg_N30;
 always @(posedge clk)
         retime_s1_32_reg_reg_N30 <= n_220;
 assign n_128 = retime_s1_32_reg_reg_N30;
 reg retime_s1_33_reg_reg_N30;
 always @(posedge clk)
         retime_s1_33_reg_reg_N30 <= n_213;
 assign n_129 = retime_s1_33_reg_reg_N30;
 reg retime_s1_34_reg_reg_N30;
 always @(posedge clk)
         retime_s1_34_reg_reg_N30 <= n_209;
 assign n_130 = retime_s1_34_reg_reg_N30;
 reg retime_s1_35_reg_reg_N30;
 always @(posedge clk)
         retime_s1_35_reg_reg_N30 <= n_203;
 assign n_131 = retime_s1_35_reg_reg_N30;
 reg retime_s1_36_reg_reg_N30;
 always @(posedge clk)
         retime_s1_36_reg_reg_N30 <= n_200;
 assign n_132 = retime_s1_36_reg_reg_N30;
 reg retime_s1_37_reg_reg_N30;
 always @(posedge clk)
         retime_s1_37_reg_reg_N30 <= n_7;
 assign n_133 = retime_s1_37_reg_reg_N30;
 reg retime_s1_38_reg_reg_N30;
 always @(posedge clk)
         retime_s1_38_reg_reg_N30 <= n_420;
 assign n_134 = retime_s1_38_reg_reg_N30;
 reg retime_s1_39_reg_reg_N30;
 always @(posedge clk)
         retime_s1_39_reg_reg_N30 <= n_0;
 assign n_135 = retime_s1_39_reg_reg_N30;
 reg retime_s1_40_reg_reg_N30;
 always @(posedge clk)
         retime_s1_40_reg_reg_N30 <= n_253;
 assign n_136 = retime_s1_40_reg_reg_N30;
 reg retime_s1_41_reg_reg_N30;
 always @(posedge clk)
         retime_s1_41_reg_reg_N30 <= n_245;
 assign n_137 = retime_s1_41_reg_reg_N30;
 reg retime_s1_42_reg_reg_N30;
 always @(posedge clk)
         retime_s1_42_reg_reg_N30 <= n_374;
 assign n_138 = retime_s1_42_reg_reg_N30;
 reg retime_s1_43_reg_reg_N30;
 always @(posedge clk)
         retime_s1_43_reg_reg_N30 <= n_18;
 assign n_139 = retime_s1_43_reg_reg_N30;
 reg retime_s1_44_reg_reg_N30;
 always @(posedge clk)
         retime_s1_44_reg_reg_N30 <= n_425;
 assign n_140 = retime_s1_44_reg_reg_N30;
 reg retime_s1_45_reg_reg_N30;
 always @(posedge clk)
         retime_s1_45_reg_reg_N30 <= n_3;
 assign n_141 = retime_s1_45_reg_reg_N30;
 reg retime_s1_46_reg_reg_N30;
 always @(posedge clk)
         retime_s1_46_reg_reg_N30 <= n_255;
 assign n_142 = retime_s1_46_reg_reg_N30;
 reg retime_s1_47_reg_reg_N30;
 always @(posedge clk)
         retime_s1_47_reg_reg_N30 <= n_247;
 assign n_143 = retime_s1_47_reg_reg_N30;
 reg retime_s1_48_reg_reg_N30;
 always @(posedge clk)
         retime_s1_48_reg_reg_N30 <= n_20;
 assign n_144 = retime_s1_48_reg_reg_N30;
 reg retime_s1_49_reg_reg_N30;
 always @(posedge clk)
         retime_s1_49_reg_reg_N30 <= n_34;
 assign n_145 = retime_s1_49_reg_reg_N30;
 reg retime_s1_50_reg_reg_N30;
 always @(posedge clk)
         retime_s1_50_reg_reg_N30 <= n_418;
 assign n_146 = retime_s1_50_reg_reg_N30;
 reg retime_s1_51_reg_reg_N30;
 always @(posedge clk)
         retime_s1_51_reg_reg_N30 <= n_423;
 assign n_147 = retime_s1_51_reg_reg_N30;
 reg retime_s1_52_reg_reg_N30;
 always @(posedge clk)
         retime_s1_52_reg_reg_N30 <= n_410;
 assign n_148 = retime_s1_52_reg_reg_N30;
 reg retime_s1_53_reg_reg_N30;
 always @(posedge clk)
         retime_s1_53_reg_reg_N30 <= n_417;
 assign n_149 = retime_s1_53_reg_reg_N30;
 reg retime_s1_54_reg_reg_N30;
 always @(posedge clk)
         retime_s1_54_reg_reg_N30 <= n_198;
 assign n_150 = retime_s1_54_reg_reg_N30;
 reg retime_s1_55_reg_reg_N30;
 always @(posedge clk)
         retime_s1_55_reg_reg_N30 <= n_227;
 assign n_151 = retime_s1_55_reg_reg_N30;
 reg retime_s1_56_reg_reg_N30;
 always @(posedge clk)
         retime_s1_56_reg_reg_N30 <= n_233;
 assign n_152 = retime_s1_56_reg_reg_N30;
 reg retime_s1_57_reg_reg_N30;
 always @(posedge clk)
         retime_s1_57_reg_reg_N30 <= n_415;
 assign n_153 = retime_s1_57_reg_reg_N30;
 reg retime_s1_58_reg_reg_N30;
 always @(posedge clk)
         retime_s1_58_reg_reg_N30 <= n_421;
 assign n_154 = retime_s1_58_reg_reg_N30;
 reg retime_s1_59_reg_reg_N30;
 always @(posedge clk)
         retime_s1_59_reg_reg_N30 <= n_411;
 assign mul_72_11_n_38 = retime_s1_59_reg_reg_N30;
 reg retime_s1_60_reg_reg_N30;
 always @(posedge clk)
         if (csa_tree_add_69_2_groupi_n_1405)
         retime_s1_60_reg_reg_N30 <= n_427;
     else
         retime_s1_60_reg_reg_N30 <= csa_tree_add_69_2_groupi_n_1420;
 assign n_155 = retime_s1_60_reg_reg_N30;
 reg retime_s1_61_reg_reg_N30;
 always @(posedge clk)
         retime_s1_61_reg_reg_N30 <= n_409;
 assign n_156 = retime_s1_61_reg_reg_N30;
 reg retime_s1_62_reg_reg_N30;
 always @(posedge clk)
         retime_s1_62_reg_reg_N30 <= n_378;
 assign n_157 = retime_s1_62_reg_reg_N30;
 reg retime_s1_63_reg_reg_N30;
 always @(posedge clk)
         retime_s1_63_reg_reg_N30 <= n_60;
 assign n_158 = retime_s1_63_reg_reg_N30;
 reg retime_s1_64_reg_reg_N30;
 always @(posedge clk)
         retime_s1_64_reg_reg_N30 <= n_61;
 assign n_159 = retime_s1_64_reg_reg_N30;
 reg retime_s1_65_reg_reg_N30;
 always @(posedge clk)
         retime_s1_65_reg_reg_N30 <= n_413;
 assign n_160 = retime_s1_65_reg_reg_N30;
 reg retime_s1_66_reg_reg_N30;
 always @(posedge clk)
         retime_s1_66_reg_reg_N30 <= n_424;
 assign n_161 = retime_s1_66_reg_reg_N30;
 reg retime_s1_67_reg_reg_N30;
 always @(posedge clk)
         retime_s1_67_reg_reg_N30 <= n_426;
 assign n_162 = retime_s1_67_reg_reg_N30;
 reg retime_s1_68_reg_reg_N30;
 always @(posedge clk)
         retime_s1_68_reg_reg_N30 <= n_422;
 assign n_163 = retime_s1_68_reg_reg_N30;
 reg retime_s1_69_reg_reg_N30;
 always @(posedge clk)
         retime_s1_69_reg_reg_N30 <= {in3[29]};
 assign n_164 = retime_s1_69_reg_reg_N30;
 reg retime_s1_70_reg_reg_N30;
 always @(posedge clk)
         retime_s1_70_reg_reg_N30 <= {in3[28]};
 assign n_165 = retime_s1_70_reg_reg_N30;
 reg retime_s1_71_reg_reg_N30;
 always @(posedge clk)
         if (csa_tree_add_69_2_groupi_n_1567)
         retime_s1_71_reg_reg_N30 <= n_428;
     else
         retime_s1_71_reg_reg_N30 <= csa_tree_add_69_2_groupi_n_1514;
 assign n_166 = retime_s1_71_reg_reg_N30;
 reg retime_s1_72_reg_reg_N30;
 always @(posedge clk)
         retime_s1_72_reg_reg_N30 <= n_219;
 assign n_167 = retime_s1_72_reg_reg_N30;
 reg retime_s1_73_reg_reg_N30;
 always @(posedge clk)
         retime_s1_73_reg_reg_N30 <= n_218;
 assign n_168 = retime_s1_73_reg_reg_N30;
 reg retime_s1_74_reg_reg_N30;
 always @(posedge clk)
         retime_s1_74_reg_reg_N30 <= n_412;
 assign n_169 = retime_s1_74_reg_reg_N30;
 reg retime_s1_75_reg_reg_N30;
 always @(posedge clk)
         retime_s1_75_reg_reg_N30 <= {in3[30]};
 assign n_170 = retime_s1_75_reg_reg_N30;
 reg retime_s1_76_reg_reg_N30;
 always @(posedge clk)
         retime_s1_76_reg_reg_N30 <= n_224;
 assign n_171 = retime_s1_76_reg_reg_N30;
 reg retime_s1_77_reg_reg_N30;
 always @(posedge clk)
         retime_s1_77_reg_reg_N30 <= n_235;
 assign n_172 = retime_s1_77_reg_reg_N30;
 assign add_59_2_n_10 = ({in8[2]} & {in9[2]});
 assign add_59_2_n_68 = ~(add_59_2_n_63 | add_59_2_n_24);
 assign n_379 = ~(add_59_2_n_9 & (add_59_2_n_18 & add_59_2_n_43));
 assign n_382 = ~add_59_2_n_64;
 assign add_59_2_n_64 = ~(add_59_2_n_60 | (add_59_2_n_56 & (add_59_2_n_21 & add_59_2_n_3)));
 assign add_59_2_n_63 = ~(add_59_2_n_58 | add_59_2_n_15);
 assign add_59_2_n_60 = ~(add_59_2_n_59 | add_59_2_n_3);
 assign add_59_2_n_59 = ~(add_59_2_n_55 | add_59_2_n_20);
 assign add_59_2_n_58 = ~(add_59_2_n_6 | add_59_2_n_38);
 assign add_59_2_n_56 = ~add_59_2_n_55;
 assign add_59_2_n_55 = ~(add_59_2_n_52 | add_59_2_n_25);
 assign add_59_2_n_52 = ~(add_59_2_n_50 | add_59_2_n_2);
 assign add_59_2_n_50 = ~(add_59_2_n_11 | add_59_2_n_28);
 assign add_59_2_n_43 = ~(add_59_2_n_7 | add_59_2_n_34);
 assign add_59_2_n_42 = ~(add_59_2_n_40 | add_59_2_n_27);
 assign add_59_2_n_40 = ~(add_59_2_n_19 | add_59_2_n_16);
 assign add_59_2_n_38 = ~(add_59_2_n_17 & (add_59_2_n_14 | add_59_2_n_21));
 assign add_59_2_n_34 = ~(add_59_2_n_22 | add_59_2_n_23);
 assign add_59_2_n_37 = ~(add_59_2_n_28 | add_59_2_n_2);
 assign add_59_2_n_36 = ~(add_59_2_n_25 | add_59_2_n_20);
 assign add_59_2_n_33 = ~(add_59_2_n_19 | add_59_2_n_27);
 assign add_59_2_n_35 = ~(add_59_2_n_15 | add_59_2_n_22);
 assign add_59_2_n_32 = ~(add_59_2_n_25 | add_59_2_n_14);
 assign add_59_2_n_31 = ~(add_59_2_n_13 | add_59_2_n_10);
 assign add_59_2_n_30 = ~(add_59_2_n_15 | add_59_2_n_24);
 assign add_59_2_n_27 = ~add_59_2_n_26;
 assign add_59_2_n_24 = ~add_59_2_n_23;
 assign add_59_2_n_20 = ~add_59_2_n_21;
 assign add_59_2_n_28 = ~({in8[3]} | {in9[3]});
 assign add_59_2_n_26 = ~({in8[1]} & {in9[1]});
 assign add_59_2_n_25 = ~({in8[4]} | {in9[4]});
 assign add_59_2_n_23 = ~({in8[6]} & {in9[6]});
 assign add_59_2_n_22 = ~({in8[7]} | {in9[7]});
 assign add_59_2_n_21 = ~({in8[4]} & {in9[4]});
 assign add_59_2_n_19 = ~({in8[1]} | {in9[1]});
 assign add_59_2_n_18 = ~({in8[7]} & {in9[7]});
 assign add_59_2_n_17 = ~({in8[5]} & {in9[5]});
 assign add_59_2_n_16 = ~({in8[0]} & {in9[0]});
 assign add_59_2_n_15 = ~({in8[6]} | {in9[6]});
 assign add_59_2_n_14 = ~({in8[5]} | {in9[5]});
 assign add_59_2_n_13 = ~({in8[2]} | {in9[2]});
 assign add_59_2_n_12 = ~(add_59_2_n_42 | add_59_2_n_13);
 assign add_59_2_n_11 = ~(add_59_2_n_12 | add_59_2_n_10);
 assign add_59_2_n_9 = ~(add_59_2_n_32 & (add_59_2_n_35 & ~add_59_2_n_52));
 assign add_59_2_n_7 = (add_59_2_n_38 & add_59_2_n_35);
 assign add_59_2_n_6 = ~(add_59_2_n_52 | ~add_59_2_n_32);
 assign add_59_2_n_5 = ~(add_59_2_n_26 & ~add_59_2_n_19);
 assign add_59_2_n_4 = ~(add_59_2_n_22 | ~add_59_2_n_18);
 assign add_59_2_n_3 = ~(add_59_2_n_14 | ~add_59_2_n_17);
 assign add_59_2_n_2 = ({in8[3]} & {in9[3]});
 assign add_63_2_n_10 = ({in5[2]} & {in6[2]});
 assign add_63_2_n_68 = ~(add_63_2_n_63 | add_63_2_n_24);
 assign n_388 = ~(add_63_2_n_9 & (add_63_2_n_18 & add_63_2_n_43));
 assign n_391 = ~add_63_2_n_64;
 assign add_63_2_n_64 = ~(add_63_2_n_60 | (add_63_2_n_56 & (add_63_2_n_21 & add_63_2_n_3)));
 assign add_63_2_n_63 = ~(add_63_2_n_58 | add_63_2_n_15);
 assign add_63_2_n_60 = ~(add_63_2_n_59 | add_63_2_n_3);
 assign add_63_2_n_59 = ~(add_63_2_n_55 | add_63_2_n_20);
 assign add_63_2_n_58 = ~(add_63_2_n_6 | add_63_2_n_38);
 assign add_63_2_n_56 = ~add_63_2_n_55;
 assign add_63_2_n_55 = ~(add_63_2_n_52 | add_63_2_n_25);
 assign add_63_2_n_52 = ~(add_63_2_n_50 | add_63_2_n_2);
 assign add_63_2_n_50 = ~(add_63_2_n_11 | add_63_2_n_28);
 assign add_63_2_n_43 = ~(add_63_2_n_7 | add_63_2_n_34);
 assign add_63_2_n_42 = ~(add_63_2_n_40 | add_63_2_n_27);
 assign add_63_2_n_40 = ~(add_63_2_n_19 | add_63_2_n_16);
 assign add_63_2_n_38 = ~(add_63_2_n_17 & (add_63_2_n_14 | add_63_2_n_21));
 assign add_63_2_n_34 = ~(add_63_2_n_22 | add_63_2_n_23);
 assign add_63_2_n_37 = ~(add_63_2_n_28 | add_63_2_n_2);
 assign add_63_2_n_36 = ~(add_63_2_n_25 | add_63_2_n_20);
 assign add_63_2_n_33 = ~(add_63_2_n_19 | add_63_2_n_27);
 assign add_63_2_n_35 = ~(add_63_2_n_15 | add_63_2_n_22);
 assign add_63_2_n_32 = ~(add_63_2_n_25 | add_63_2_n_14);
 assign add_63_2_n_31 = ~(add_63_2_n_13 | add_63_2_n_10);
 assign add_63_2_n_30 = ~(add_63_2_n_15 | add_63_2_n_24);
 assign add_63_2_n_27 = ~add_63_2_n_26;
 assign add_63_2_n_24 = ~add_63_2_n_23;
 assign add_63_2_n_20 = ~add_63_2_n_21;
 assign add_63_2_n_28 = ~({in5[3]} | {in6[3]});
 assign add_63_2_n_26 = ~({in5[1]} & {in6[1]});
 assign add_63_2_n_25 = ~({in5[4]} | {in6[4]});
 assign add_63_2_n_23 = ~({in5[6]} & {in6[6]});
 assign add_63_2_n_22 = ~({in5[7]} | {in6[7]});
 assign add_63_2_n_21 = ~({in5[4]} & {in6[4]});
 assign add_63_2_n_19 = ~({in5[1]} | {in6[1]});
 assign add_63_2_n_18 = ~({in5[7]} & {in6[7]});
 assign add_63_2_n_17 = ~({in5[5]} & {in6[5]});
 assign add_63_2_n_16 = ~({in5[0]} & {in6[0]});
 assign add_63_2_n_15 = ~({in5[6]} | {in6[6]});
 assign add_63_2_n_14 = ~({in5[5]} | {in6[5]});
 assign add_63_2_n_13 = ~({in5[2]} | {in6[2]});
 assign add_63_2_n_12 = ~(add_63_2_n_42 | add_63_2_n_13);
 assign add_63_2_n_11 = ~(add_63_2_n_12 | add_63_2_n_10);
 assign add_63_2_n_9 = ~(add_63_2_n_32 & (add_63_2_n_35 & ~add_63_2_n_52));
 assign add_63_2_n_7 = (add_63_2_n_38 & add_63_2_n_35);
 assign add_63_2_n_6 = ~(add_63_2_n_52 | ~add_63_2_n_32);
 assign add_63_2_n_5 = ~(add_63_2_n_26 & ~add_63_2_n_19);
 assign add_63_2_n_4 = ~(add_63_2_n_22 | ~add_63_2_n_18);
 assign add_63_2_n_3 = ~(add_63_2_n_14 | ~add_63_2_n_17);
 assign add_63_2_n_2 = ({in5[3]} & {in6[3]});
 assign csa_tree_add_55_2_groupi_n_228 = ~({in3[26]} & ~csa_tree_add_55_2_groupi_n_226);
 assign csa_tree_add_55_2_groupi_n_226 = ~({in3[25]} & ~csa_tree_add_55_2_groupi_n_224);
 assign csa_tree_add_55_2_groupi_n_224 = ~({in3[24]} & ~csa_tree_add_55_2_groupi_n_222);
 assign csa_tree_add_55_2_groupi_n_222 = ~({in3[23]} & ~csa_tree_add_55_2_groupi_n_220);
 assign csa_tree_add_55_2_groupi_n_220 = ~({in3[22]} & ~csa_tree_add_55_2_groupi_n_218);
 assign csa_tree_add_55_2_groupi_n_218 = ~({in3[21]} & ~csa_tree_add_55_2_groupi_n_216);
 assign csa_tree_add_55_2_groupi_n_216 = ~({in3[20]} & ~csa_tree_add_55_2_groupi_n_214);
 assign csa_tree_add_55_2_groupi_n_214 = ~({in3[19]} & ~csa_tree_add_55_2_groupi_n_212);
 assign csa_tree_add_55_2_groupi_n_212 = ~({in3[18]} & ~csa_tree_add_55_2_groupi_n_210);
 assign csa_tree_add_55_2_groupi_n_210 = ~({in3[17]} & ~csa_tree_add_55_2_groupi_n_208);
 assign csa_tree_add_55_2_groupi_n_208 = ~(csa_tree_add_55_2_groupi_n_207 & {in3[16]});
 assign csa_tree_add_55_2_groupi_n_186 = ((csa_tree_add_55_2_groupi_n_162 & csa_tree_add_55_2_groupi_n_165)
    | ((csa_tree_add_55_2_groupi_n_165 & csa_tree_add_55_2_groupi_n_147) | (csa_tree_add_55_2_groupi_n_147
    & csa_tree_add_55_2_groupi_n_162)));
 assign csa_tree_add_55_2_groupi_n_187 = (csa_tree_add_55_2_groupi_n_165 ^ (csa_tree_add_55_2_groupi_n_147
    ^ csa_tree_add_55_2_groupi_n_162));
 assign csa_tree_add_55_2_groupi_n_184 = ((csa_tree_add_55_2_groupi_n_164 & csa_tree_add_55_2_groupi_n_169)
    | ((csa_tree_add_55_2_groupi_n_169 & csa_tree_add_55_2_groupi_n_151) | (csa_tree_add_55_2_groupi_n_151
    & csa_tree_add_55_2_groupi_n_164)));
 assign csa_tree_add_55_2_groupi_n_185 = (csa_tree_add_55_2_groupi_n_169 ^ (csa_tree_add_55_2_groupi_n_151
    ^ csa_tree_add_55_2_groupi_n_164));
 assign csa_tree_add_55_2_groupi_n_180 = ((csa_tree_add_55_2_groupi_n_158 & csa_tree_add_55_2_groupi_n_163)
    | ((csa_tree_add_55_2_groupi_n_163 & csa_tree_add_55_2_groupi_n_145) | (csa_tree_add_55_2_groupi_n_145
    & csa_tree_add_55_2_groupi_n_158)));
 assign csa_tree_add_55_2_groupi_n_181 = (csa_tree_add_55_2_groupi_n_163 ^ (csa_tree_add_55_2_groupi_n_145
    ^ csa_tree_add_55_2_groupi_n_158));
 assign csa_tree_add_55_2_groupi_n_178 = ((csa_tree_add_55_2_groupi_n_159 & csa_tree_add_55_2_groupi_n_154)
    | ((csa_tree_add_55_2_groupi_n_154 & csa_tree_add_55_2_groupi_n_149) | (csa_tree_add_55_2_groupi_n_149
    & csa_tree_add_55_2_groupi_n_159)));
 assign csa_tree_add_55_2_groupi_n_179 = (csa_tree_add_55_2_groupi_n_154 ^ (csa_tree_add_55_2_groupi_n_149
    ^ csa_tree_add_55_2_groupi_n_159));
 assign csa_tree_add_55_2_groupi_n_174 = ((csa_tree_add_55_2_groupi_n_168 & csa_tree_add_55_2_groupi_n_150)
    | ((csa_tree_add_55_2_groupi_n_150 & csa_tree_add_55_2_groupi_n_141) | (csa_tree_add_55_2_groupi_n_141
    & csa_tree_add_55_2_groupi_n_168)));
 assign csa_tree_add_55_2_groupi_n_175 = (csa_tree_add_55_2_groupi_n_150 ^ (csa_tree_add_55_2_groupi_n_141
    ^ csa_tree_add_55_2_groupi_n_168));
 assign csa_tree_add_55_2_groupi_n_172 = ((csa_tree_add_55_2_groupi_n_140 & csa_tree_add_55_2_groupi_n_124)
    | ((csa_tree_add_55_2_groupi_n_124 & csa_tree_add_55_2_groupi_n_137) | (csa_tree_add_55_2_groupi_n_137
    & csa_tree_add_55_2_groupi_n_140)));
 assign csa_tree_add_55_2_groupi_n_173 = (csa_tree_add_55_2_groupi_n_124 ^ (csa_tree_add_55_2_groupi_n_137
    ^ csa_tree_add_55_2_groupi_n_140));
 assign csa_tree_add_55_2_groupi_n_170 = ((csa_tree_add_55_2_groupi_n_155 & csa_tree_add_55_2_groupi_n_142)
    | ((csa_tree_add_55_2_groupi_n_142 & csa_tree_add_55_2_groupi_n_135) | (csa_tree_add_55_2_groupi_n_135
    & csa_tree_add_55_2_groupi_n_155)));
 assign csa_tree_add_55_2_groupi_n_171 = (csa_tree_add_55_2_groupi_n_142 ^ (csa_tree_add_55_2_groupi_n_135
    ^ csa_tree_add_55_2_groupi_n_155));
 assign csa_tree_add_55_2_groupi_n_168 = ((csa_tree_add_55_2_groupi_n_146 & csa_tree_add_55_2_groupi_n_91)
    | ((csa_tree_add_55_2_groupi_n_91 & csa_tree_add_55_2_groupi_n_132) | (csa_tree_add_55_2_groupi_n_132
    & csa_tree_add_55_2_groupi_n_146)));
 assign csa_tree_add_55_2_groupi_n_169 = (csa_tree_add_55_2_groupi_n_91 ^ (csa_tree_add_55_2_groupi_n_132
    ^ csa_tree_add_55_2_groupi_n_146));
 assign csa_tree_add_55_2_groupi_n_164 = ((csa_tree_add_55_2_groupi_n_144 & csa_tree_add_55_2_groupi_n_128)
    | ((csa_tree_add_55_2_groupi_n_128 & csa_tree_add_55_2_groupi_n_133) | (csa_tree_add_55_2_groupi_n_133
    & csa_tree_add_55_2_groupi_n_144)));
 assign csa_tree_add_55_2_groupi_n_165 = (csa_tree_add_55_2_groupi_n_128 ^ (csa_tree_add_55_2_groupi_n_133
    ^ csa_tree_add_55_2_groupi_n_144));
 assign csa_tree_add_55_2_groupi_n_162 = ((csa_tree_add_55_2_groupi_n_148 & csa_tree_add_55_2_groupi_n_118)
    | ((csa_tree_add_55_2_groupi_n_118 & csa_tree_add_55_2_groupi_n_129) | (csa_tree_add_55_2_groupi_n_129
    & csa_tree_add_55_2_groupi_n_148)));
 assign csa_tree_add_55_2_groupi_n_163 = (csa_tree_add_55_2_groupi_n_118 ^ (csa_tree_add_55_2_groupi_n_129
    ^ csa_tree_add_55_2_groupi_n_148));
 assign csa_tree_add_55_2_groupi_n_160 = ((csa_tree_add_55_2_groupi_n_136 & csa_tree_add_55_2_groupi_n_86)
    | ((csa_tree_add_55_2_groupi_n_86 & csa_tree_add_55_2_groupi_n_89) | (csa_tree_add_55_2_groupi_n_89 &
    csa_tree_add_55_2_groupi_n_136)));
 assign csa_tree_add_55_2_groupi_n_161 = (csa_tree_add_55_2_groupi_n_86 ^ (csa_tree_add_55_2_groupi_n_89
    ^ csa_tree_add_55_2_groupi_n_136));
 assign csa_tree_add_55_2_groupi_n_158 = ((csa_tree_add_55_2_groupi_n_134 & csa_tree_add_55_2_groupi_n_119)
    | ((csa_tree_add_55_2_groupi_n_119 & csa_tree_add_55_2_groupi_n_113) | (csa_tree_add_55_2_groupi_n_113
    & csa_tree_add_55_2_groupi_n_134)));
 assign csa_tree_add_55_2_groupi_n_159 = (csa_tree_add_55_2_groupi_n_119 ^ (csa_tree_add_55_2_groupi_n_113
    ^ csa_tree_add_55_2_groupi_n_134));
 assign csa_tree_add_55_2_groupi_n_156 = ((csa_tree_add_55_2_groupi_n_143 & csa_tree_add_55_2_groupi_n_120)
    | ((csa_tree_add_55_2_groupi_n_120 & csa_tree_add_55_2_groupi_n_105) | (csa_tree_add_55_2_groupi_n_105
    & csa_tree_add_55_2_groupi_n_143)));
 assign csa_tree_add_55_2_groupi_n_157 = (csa_tree_add_55_2_groupi_n_120 ^ (csa_tree_add_55_2_groupi_n_105
    ^ csa_tree_add_55_2_groupi_n_143));
 assign csa_tree_add_55_2_groupi_n_154 = ((csa_tree_add_55_2_groupi_n_104 & csa_tree_add_55_2_groupi_n_101)
    | ((csa_tree_add_55_2_groupi_n_101 & csa_tree_add_55_2_groupi_n_103) | (csa_tree_add_55_2_groupi_n_103
    & csa_tree_add_55_2_groupi_n_104)));
 assign csa_tree_add_55_2_groupi_n_155 = (csa_tree_add_55_2_groupi_n_101 ^ (csa_tree_add_55_2_groupi_n_103
    ^ csa_tree_add_55_2_groupi_n_104));
 assign csa_tree_add_55_2_groupi_n_150 = ((csa_tree_add_55_2_groupi_n_85 & csa_tree_add_55_2_groupi_n_110)
    | ((csa_tree_add_55_2_groupi_n_110 & csa_tree_add_55_2_groupi_n_106) | (csa_tree_add_55_2_groupi_n_106
    & csa_tree_add_55_2_groupi_n_85)));
 assign csa_tree_add_55_2_groupi_n_151 = (csa_tree_add_55_2_groupi_n_110 ^ (csa_tree_add_55_2_groupi_n_106
    ^ csa_tree_add_55_2_groupi_n_85));
 assign csa_tree_add_55_2_groupi_n_148 = ((csa_tree_add_55_2_groupi_n_109 & csa_tree_add_55_2_groupi_n_102)
    | ((csa_tree_add_55_2_groupi_n_102 & csa_tree_add_55_2_groupi_n_100) | (csa_tree_add_55_2_groupi_n_100
    & csa_tree_add_55_2_groupi_n_109)));
 assign csa_tree_add_55_2_groupi_n_149 = (csa_tree_add_55_2_groupi_n_102 ^ (csa_tree_add_55_2_groupi_n_100
    ^ csa_tree_add_55_2_groupi_n_109));
 assign csa_tree_add_55_2_groupi_n_146 = ((csa_tree_add_55_2_groupi_n_107 & csa_tree_add_55_2_groupi_n_92)
    | ((csa_tree_add_55_2_groupi_n_92 & csa_tree_add_55_2_groupi_n_111) | (csa_tree_add_55_2_groupi_n_111
    & csa_tree_add_55_2_groupi_n_107)));
 assign csa_tree_add_55_2_groupi_n_147 = (csa_tree_add_55_2_groupi_n_92 ^ (csa_tree_add_55_2_groupi_n_111
    ^ csa_tree_add_55_2_groupi_n_107));
 assign csa_tree_add_55_2_groupi_n_144 = ((csa_tree_add_55_2_groupi_n_93 & csa_tree_add_55_2_groupi_n_108)
    | ((csa_tree_add_55_2_groupi_n_108 & csa_tree_add_55_2_groupi_n_99) | (csa_tree_add_55_2_groupi_n_99
    & csa_tree_add_55_2_groupi_n_93)));
 assign csa_tree_add_55_2_groupi_n_145 = (csa_tree_add_55_2_groupi_n_108 ^ (csa_tree_add_55_2_groupi_n_99
    ^ csa_tree_add_55_2_groupi_n_93));
 assign csa_tree_add_55_2_groupi_n_142 = ((csa_tree_add_55_2_groupi_n_117 & csa_tree_add_55_2_groupi_n_67)
    | ((csa_tree_add_55_2_groupi_n_67 & csa_tree_add_55_2_groupi_n_82) | (csa_tree_add_55_2_groupi_n_82 &
    csa_tree_add_55_2_groupi_n_117)));
 assign csa_tree_add_55_2_groupi_n_143 = (csa_tree_add_55_2_groupi_n_67 ^ (csa_tree_add_55_2_groupi_n_82
    ^ csa_tree_add_55_2_groupi_n_117));
 assign csa_tree_add_55_2_groupi_n_140 = ((csa_tree_add_55_2_groupi_n_125 & csa_tree_add_55_2_groupi_n_84)
    | ((csa_tree_add_55_2_groupi_n_84 & csa_tree_add_55_2_groupi_n_97) | (csa_tree_add_55_2_groupi_n_97 &
    csa_tree_add_55_2_groupi_n_125)));
 assign csa_tree_add_55_2_groupi_n_141 = (csa_tree_add_55_2_groupi_n_84 ^ (csa_tree_add_55_2_groupi_n_97
    ^ csa_tree_add_55_2_groupi_n_125));
 assign csa_tree_add_55_2_groupi_n_138 = ((csa_tree_add_55_2_groupi_n_121 & csa_tree_add_55_2_groupi_n_94)
    | ((csa_tree_add_55_2_groupi_n_94 & csa_tree_add_55_2_groupi_n_83) | (csa_tree_add_55_2_groupi_n_83 &
    csa_tree_add_55_2_groupi_n_121)));
 assign csa_tree_add_55_2_groupi_n_139 = (csa_tree_add_55_2_groupi_n_94 ^ (csa_tree_add_55_2_groupi_n_83
    ^ csa_tree_add_55_2_groupi_n_121));
 assign csa_tree_add_55_2_groupi_n_136 = ((csa_tree_add_55_2_groupi_n_87 & csa_tree_add_55_2_groupi_n_44)
    | ((csa_tree_add_55_2_groupi_n_44 & csa_tree_add_55_2_groupi_n_96) | (csa_tree_add_55_2_groupi_n_96 &
    csa_tree_add_55_2_groupi_n_87)));
 assign csa_tree_add_55_2_groupi_n_137 = (csa_tree_add_55_2_groupi_n_44 ^ (csa_tree_add_55_2_groupi_n_96
    ^ csa_tree_add_55_2_groupi_n_87));
 assign csa_tree_add_55_2_groupi_n_134 = ((csa_tree_add_55_2_groupi_n_116 & csa_tree_add_55_2_groupi_n_66)
    | ((csa_tree_add_55_2_groupi_n_66 & csa_tree_add_55_2_groupi_n_69) | (csa_tree_add_55_2_groupi_n_69 &
    csa_tree_add_55_2_groupi_n_116)));
 assign csa_tree_add_55_2_groupi_n_135 = (csa_tree_add_55_2_groupi_n_66 ^ (csa_tree_add_55_2_groupi_n_69
    ^ csa_tree_add_55_2_groupi_n_116));
 assign csa_tree_add_55_2_groupi_n_132 = ((csa_tree_add_55_2_groupi_n_98 & csa_tree_add_55_2_groupi_n_46)
    | ((csa_tree_add_55_2_groupi_n_46 & csa_tree_add_55_2_groupi_n_80) | (csa_tree_add_55_2_groupi_n_80 &
    csa_tree_add_55_2_groupi_n_98)));
 assign csa_tree_add_55_2_groupi_n_133 = (csa_tree_add_55_2_groupi_n_46 ^ (csa_tree_add_55_2_groupi_n_80
    ^ csa_tree_add_55_2_groupi_n_98));
 assign csa_tree_add_55_2_groupi_n_130 = ((csa_tree_add_55_2_groupi_n_95 & csa_tree_add_55_2_groupi_n_64)
    | ((csa_tree_add_55_2_groupi_n_64 & csa_tree_add_55_2_groupi_n_73) | (csa_tree_add_55_2_groupi_n_73 &
    csa_tree_add_55_2_groupi_n_95)));
 assign csa_tree_add_55_2_groupi_n_131 = (csa_tree_add_55_2_groupi_n_64 ^ (csa_tree_add_55_2_groupi_n_73
    ^ csa_tree_add_55_2_groupi_n_95));
 assign csa_tree_add_55_2_groupi_n_128 = ((csa_tree_add_55_2_groupi_n_112 & csa_tree_add_55_2_groupi_n_70)
    | ((csa_tree_add_55_2_groupi_n_70 & csa_tree_add_55_2_groupi_n_81) | (csa_tree_add_55_2_groupi_n_81 &
    csa_tree_add_55_2_groupi_n_112)));
 assign csa_tree_add_55_2_groupi_n_129 = (csa_tree_add_55_2_groupi_n_70 ^ (csa_tree_add_55_2_groupi_n_81
    ^ csa_tree_add_55_2_groupi_n_112));
 assign csa_tree_add_55_2_groupi_n_124 = ((csa_tree_add_55_2_groupi_n_90 & csa_tree_add_55_2_groupi_n_11)
    | ((csa_tree_add_55_2_groupi_n_11 & csa_tree_add_55_2_groupi_n_47) | (csa_tree_add_55_2_groupi_n_47 &
    csa_tree_add_55_2_groupi_n_90)));
 assign csa_tree_add_55_2_groupi_n_125 = (csa_tree_add_55_2_groupi_n_11 ^ (csa_tree_add_55_2_groupi_n_47
    ^ csa_tree_add_55_2_groupi_n_90));
 assign csa_tree_add_55_2_groupi_n_122 = ((csa_tree_add_55_2_groupi_n_88 & csa_tree_add_55_2_groupi_n_9)
    | ((csa_tree_add_55_2_groupi_n_9 & {in3[14]}) | ({in3[14]} & csa_tree_add_55_2_groupi_n_88)));
 assign csa_tree_add_55_2_groupi_n_123 = (csa_tree_add_55_2_groupi_n_9 ^ ({in3[14]} ^ csa_tree_add_55_2_groupi_n_88));
 assign csa_tree_add_55_2_groupi_n_120 = ((csa_tree_add_55_2_groupi_n_77 & csa_tree_add_55_2_groupi_n_4)
    | ((csa_tree_add_55_2_groupi_n_4 & csa_tree_add_55_2_groupi_n_72) | (csa_tree_add_55_2_groupi_n_72 &
    csa_tree_add_55_2_groupi_n_77)));
 assign csa_tree_add_55_2_groupi_n_121 = (csa_tree_add_55_2_groupi_n_4 ^ (csa_tree_add_55_2_groupi_n_72
    ^ csa_tree_add_55_2_groupi_n_77));
 assign csa_tree_add_55_2_groupi_n_118 = ((csa_tree_add_55_2_groupi_n_71 & csa_tree_add_55_2_groupi_n_50)
    | ((csa_tree_add_55_2_groupi_n_50 & csa_tree_add_55_2_groupi_n_68) | (csa_tree_add_55_2_groupi_n_68 &
    csa_tree_add_55_2_groupi_n_71)));
 assign csa_tree_add_55_2_groupi_n_119 = (csa_tree_add_55_2_groupi_n_50 ^ (csa_tree_add_55_2_groupi_n_68
    ^ csa_tree_add_55_2_groupi_n_71));
 assign csa_tree_add_55_2_groupi_n_116 = ((csa_tree_add_55_2_groupi_n_25 & csa_tree_add_55_2_groupi_n_7)
    | ((csa_tree_add_55_2_groupi_n_7 & csa_tree_add_55_2_groupi_n_12) | (csa_tree_add_55_2_groupi_n_12 &
    csa_tree_add_55_2_groupi_n_25)));
 assign csa_tree_add_55_2_groupi_n_117 = (csa_tree_add_55_2_groupi_n_7 ^ (csa_tree_add_55_2_groupi_n_12
    ^ csa_tree_add_55_2_groupi_n_25));
 assign csa_tree_add_55_2_groupi_n_114 = ((csa_tree_add_55_2_groupi_n_65 & csa_tree_add_55_2_groupi_n_6)
    | ((csa_tree_add_55_2_groupi_n_6 & csa_tree_add_55_2_groupi_n_52) | (csa_tree_add_55_2_groupi_n_52 &
    csa_tree_add_55_2_groupi_n_65)));
 assign csa_tree_add_55_2_groupi_n_115 = (csa_tree_add_55_2_groupi_n_6 ^ (csa_tree_add_55_2_groupi_n_52
    ^ csa_tree_add_55_2_groupi_n_65));
 assign csa_tree_add_55_2_groupi_n_112 = ((csa_tree_add_55_2_groupi_n_24 & csa_tree_add_55_2_groupi_n_48)
    | ((csa_tree_add_55_2_groupi_n_48 & csa_tree_add_55_2_groupi_n_42) | (csa_tree_add_55_2_groupi_n_42 &
    csa_tree_add_55_2_groupi_n_24)));
 assign csa_tree_add_55_2_groupi_n_113 = (csa_tree_add_55_2_groupi_n_48 ^ (csa_tree_add_55_2_groupi_n_42
    ^ csa_tree_add_55_2_groupi_n_24));
 assign csa_tree_add_55_2_groupi_n_110 = ((csa_tree_add_55_2_groupi_n_59 & csa_tree_add_55_2_groupi_n_2)
    | ((csa_tree_add_55_2_groupi_n_2 & {in3[9]}) | ({in3[9]} & csa_tree_add_55_2_groupi_n_59)));
 assign csa_tree_add_55_2_groupi_n_111 = (csa_tree_add_55_2_groupi_n_2 ^ ({in3[9]} ^ csa_tree_add_55_2_groupi_n_59));
 assign csa_tree_add_55_2_groupi_n_108 = ((csa_tree_add_55_2_groupi_n_22 & csa_tree_add_55_2_groupi_n_5)
    | ((csa_tree_add_55_2_groupi_n_5 & csa_tree_add_55_2_groupi_n_34) | (csa_tree_add_55_2_groupi_n_34 &
    csa_tree_add_55_2_groupi_n_22)));
 assign csa_tree_add_55_2_groupi_n_109 = (csa_tree_add_55_2_groupi_n_5 ^ (csa_tree_add_55_2_groupi_n_34
    ^ csa_tree_add_55_2_groupi_n_22));
 assign csa_tree_add_55_2_groupi_n_106 = ((csa_tree_add_55_2_groupi_n_18 & csa_tree_add_55_2_groupi_n_15)
    | ((csa_tree_add_55_2_groupi_n_15 & csa_tree_add_55_2_groupi_n_8) | (csa_tree_add_55_2_groupi_n_8 & csa_tree_add_55_2_groupi_n_18)));
 assign csa_tree_add_55_2_groupi_n_107 = (csa_tree_add_55_2_groupi_n_15 ^ (csa_tree_add_55_2_groupi_n_8
    ^ csa_tree_add_55_2_groupi_n_18));
 assign csa_tree_add_55_2_groupi_n_104 = ((csa_tree_add_55_2_groupi_n_76 & csa_tree_add_55_2_groupi_n_14)
    | ((csa_tree_add_55_2_groupi_n_14 & csa_tree_add_55_2_groupi_n_10) | (csa_tree_add_55_2_groupi_n_10 &
    csa_tree_add_55_2_groupi_n_76)));
 assign csa_tree_add_55_2_groupi_n_105 = (csa_tree_add_55_2_groupi_n_14 ^ (csa_tree_add_55_2_groupi_n_10
    ^ csa_tree_add_55_2_groupi_n_76));
 assign csa_tree_add_55_2_groupi_n_102 = ((csa_tree_add_55_2_groupi_n_19 & csa_tree_add_55_2_groupi_n_51)
    | ((csa_tree_add_55_2_groupi_n_51 & csa_tree_add_55_2_groupi_n_38) | (csa_tree_add_55_2_groupi_n_38 &
    csa_tree_add_55_2_groupi_n_19)));
 assign csa_tree_add_55_2_groupi_n_103 = (csa_tree_add_55_2_groupi_n_51 ^ (csa_tree_add_55_2_groupi_n_38
    ^ csa_tree_add_55_2_groupi_n_19));
 assign csa_tree_add_55_2_groupi_n_100 = ((csa_tree_add_55_2_groupi_n_27 & csa_tree_add_55_2_groupi_n_41)
    | ((csa_tree_add_55_2_groupi_n_41 & csa_tree_add_55_2_groupi_n_13) | (csa_tree_add_55_2_groupi_n_13 &
    csa_tree_add_55_2_groupi_n_27)));
 assign csa_tree_add_55_2_groupi_n_101 = (csa_tree_add_55_2_groupi_n_41 ^ (csa_tree_add_55_2_groupi_n_13
    ^ csa_tree_add_55_2_groupi_n_27));
 assign csa_tree_add_55_2_groupi_n_98 = ((csa_tree_add_55_2_groupi_n_53 & csa_tree_add_55_2_groupi_n_0)
    | ((csa_tree_add_55_2_groupi_n_0 & csa_tree_add_55_2_groupi_n_45) | (csa_tree_add_55_2_groupi_n_45 &
    csa_tree_add_55_2_groupi_n_53)));
 assign csa_tree_add_55_2_groupi_n_99 = (csa_tree_add_55_2_groupi_n_0 ^ (csa_tree_add_55_2_groupi_n_45
    ^ csa_tree_add_55_2_groupi_n_53));
 assign csa_tree_add_55_2_groupi_n_96 = ((csa_tree_add_55_2_groupi_n_62 & csa_tree_add_55_2_groupi_n_16)
    | ((csa_tree_add_55_2_groupi_n_16 & {in3[11]}) | ({in3[11]} & csa_tree_add_55_2_groupi_n_62)));
 assign csa_tree_add_55_2_groupi_n_97 = (csa_tree_add_55_2_groupi_n_16 ^ ({in3[11]} ^ csa_tree_add_55_2_groupi_n_62));
 assign csa_tree_add_55_2_groupi_n_94 = ((csa_tree_add_55_2_groupi_n_61 & csa_tree_add_55_2_groupi_n_39)
    | ((csa_tree_add_55_2_groupi_n_39 & csa_tree_add_55_2_groupi_n_17) | (csa_tree_add_55_2_groupi_n_17 &
    csa_tree_add_55_2_groupi_n_61)));
 assign csa_tree_add_55_2_groupi_n_95 = (csa_tree_add_55_2_groupi_n_39 ^ (csa_tree_add_55_2_groupi_n_17
    ^ csa_tree_add_55_2_groupi_n_61));
 assign csa_tree_add_55_2_groupi_n_92 = ((csa_tree_add_55_2_groupi_n_21 & csa_tree_add_55_2_groupi_n_37)
    | ((csa_tree_add_55_2_groupi_n_37 & csa_tree_add_55_2_groupi_n_33) | (csa_tree_add_55_2_groupi_n_33 &
    csa_tree_add_55_2_groupi_n_21)));
 assign csa_tree_add_55_2_groupi_n_93 = (csa_tree_add_55_2_groupi_n_37 ^ (csa_tree_add_55_2_groupi_n_33
    ^ csa_tree_add_55_2_groupi_n_21));
 assign csa_tree_add_55_2_groupi_n_90 = ((csa_tree_add_55_2_groupi_n_20 & csa_tree_add_55_2_groupi_n_1)
    | ((csa_tree_add_55_2_groupi_n_1 & csa_tree_add_55_2_groupi_n_40) | (csa_tree_add_55_2_groupi_n_40 &
    csa_tree_add_55_2_groupi_n_20)));
 assign csa_tree_add_55_2_groupi_n_91 = (csa_tree_add_55_2_groupi_n_1 ^ (csa_tree_add_55_2_groupi_n_40
    ^ csa_tree_add_55_2_groupi_n_20));
 assign csa_tree_add_55_2_groupi_n_88 = ((csa_tree_add_55_2_groupi_n_30 & {in3[13]}) | (({in3[13]} &
    csa_tree_add_55_2_groupi_n_36) | (csa_tree_add_55_2_groupi_n_36 & csa_tree_add_55_2_groupi_n_30)));
 assign csa_tree_add_55_2_groupi_n_89 = ({in3[13]} ^ (csa_tree_add_55_2_groupi_n_36 ^ csa_tree_add_55_2_groupi_n_30));
 assign csa_tree_add_55_2_groupi_n_86 = ((csa_tree_add_55_2_groupi_n_29 & csa_tree_add_55_2_groupi_n_35)
    | ((csa_tree_add_55_2_groupi_n_35 & {in3[12]}) | ({in3[12]} & csa_tree_add_55_2_groupi_n_29)));
 assign csa_tree_add_55_2_groupi_n_87 = (csa_tree_add_55_2_groupi_n_35 ^ ({in3[12]} ^ csa_tree_add_55_2_groupi_n_29));
 assign csa_tree_add_55_2_groupi_n_84 = ((csa_tree_add_55_2_groupi_n_56 & csa_tree_add_55_2_groupi_n_32)
    | ((csa_tree_add_55_2_groupi_n_32 & {in3[10]}) | ({in3[10]} & csa_tree_add_55_2_groupi_n_56)));
 assign csa_tree_add_55_2_groupi_n_85 = (csa_tree_add_55_2_groupi_n_32 ^ ({in3[10]} ^ csa_tree_add_55_2_groupi_n_56));
 assign csa_tree_add_55_2_groupi_n_82 = ((csa_tree_add_55_2_groupi_n_26 & csa_tree_add_55_2_groupi_n_49)
    | ((csa_tree_add_55_2_groupi_n_49 & csa_tree_add_55_2_groupi_n_3) | (csa_tree_add_55_2_groupi_n_3 & csa_tree_add_55_2_groupi_n_26)));
 assign csa_tree_add_55_2_groupi_n_83 = (csa_tree_add_55_2_groupi_n_49 ^ (csa_tree_add_55_2_groupi_n_3
    ^ csa_tree_add_55_2_groupi_n_26));
 assign csa_tree_add_55_2_groupi_n_80 = (csa_tree_add_55_2_groupi_n_55 & {in3[8]});
 assign csa_tree_add_55_2_groupi_n_81 = (csa_tree_add_55_2_groupi_n_55 ^ {in3[8]});
 assign csa_tree_add_55_2_groupi_n_76 = (csa_tree_add_55_2_groupi_n_54 & {in3[4]});
 assign csa_tree_add_55_2_groupi_n_77 = (csa_tree_add_55_2_groupi_n_54 ^ {in3[4]});
 assign csa_tree_add_55_2_groupi_n_74 = (csa_tree_add_55_2_groupi_n_23 & {in3[1]});
 assign csa_tree_add_55_2_groupi_n_75 = (csa_tree_add_55_2_groupi_n_23 ^ {in3[1]});
 assign csa_tree_add_55_2_groupi_n_72 = (csa_tree_add_55_2_groupi_n_63 & {in3[3]});
 assign csa_tree_add_55_2_groupi_n_73 = (csa_tree_add_55_2_groupi_n_63 ^ {in3[3]});
 assign csa_tree_add_55_2_groupi_n_70 = (csa_tree_add_55_2_groupi_n_60 & {in3[7]});
 assign csa_tree_add_55_2_groupi_n_71 = (csa_tree_add_55_2_groupi_n_60 ^ {in3[7]});
 assign csa_tree_add_55_2_groupi_n_68 = (csa_tree_add_55_2_groupi_n_28 & {in3[6]});
 assign csa_tree_add_55_2_groupi_n_69 = (csa_tree_add_55_2_groupi_n_28 ^ {in3[6]});
 assign csa_tree_add_55_2_groupi_n_66 = (csa_tree_add_55_2_groupi_n_58 & {in3[5]});
 assign csa_tree_add_55_2_groupi_n_67 = (csa_tree_add_55_2_groupi_n_58 ^ {in3[5]});
 assign csa_tree_add_55_2_groupi_n_64 = (csa_tree_add_55_2_groupi_n_57 & {in3[2]});
 assign csa_tree_add_55_2_groupi_n_65 = (csa_tree_add_55_2_groupi_n_57 ^ {in3[2]});
 assign csa_tree_add_55_2_groupi_n_63 = ({in2[0]} & {in1[3]});
 assign csa_tree_add_55_2_groupi_n_62 = ({in2[4]} & {in1[7]});
 assign csa_tree_add_55_2_groupi_n_61 = ({in2[3]} & {in1[0]});
 assign csa_tree_add_55_2_groupi_n_60 = ({in2[0]} & {in1[7]});
 assign csa_tree_add_55_2_groupi_n_59 = ({in2[4]} & {in1[5]});
 assign csa_tree_add_55_2_groupi_n_58 = ({in2[0]} & {in1[5]});
 assign csa_tree_add_55_2_groupi_n_57 = ({in2[0]} & {in1[2]});
 assign csa_tree_add_55_2_groupi_n_56 = ({in2[3]} & {in1[7]});
 assign csa_tree_add_55_2_groupi_n_55 = ({in2[1]} & {in1[7]});
 assign csa_tree_add_55_2_groupi_n_54 = ({in2[0]} & {in1[4]});
 assign csa_tree_add_55_2_groupi_n_53 = ({in2[4]} & {in1[4]});
 assign csa_tree_add_55_2_groupi_n_52 = ({in2[1]} & {in1[1]});
 assign csa_tree_add_55_2_groupi_n_51 = ({in2[6]} & {in1[0]});
 assign csa_tree_add_55_2_groupi_n_50 = ({in2[5]} & {in1[2]});
 assign csa_tree_add_55_2_groupi_n_49 = ({in2[2]} & {in1[2]});
 assign csa_tree_add_55_2_groupi_n_48 = ({in2[6]} & {in1[1]});
 assign csa_tree_add_55_2_groupi_n_47 = ({in2[5]} & {in1[6]});
 assign csa_tree_add_55_2_groupi_n_46 = ({in2[7]} & {in1[2]});
 assign csa_tree_add_55_2_groupi_n_45 = ({in2[3]} & {in1[5]});
 assign csa_tree_add_55_2_groupi_n_44 = ({in2[6]} & {in1[6]});
 assign csa_tree_add_55_2_groupi_n_43 = ({in2[0]} & {in1[1]});
 assign csa_tree_add_55_2_groupi_n_42 = ({in2[2]} & {in1[5]});
 assign csa_tree_add_55_2_groupi_n_41 = ({in2[4]} & {in1[2]});
 assign csa_tree_add_55_2_groupi_n_40 = ({in2[6]} & {in1[4]});
 assign csa_tree_add_55_2_groupi_n_39 = ({in2[2]} & {in1[1]});
 assign csa_tree_add_55_2_groupi_n_38 = ({in2[2]} & {in1[4]});
 assign csa_tree_add_55_2_groupi_n_37 = ({in2[6]} & {in1[2]});
 assign csa_tree_add_55_2_groupi_n_36 = ({in2[7]} & {in1[6]});
 assign csa_tree_add_55_2_groupi_n_35 = ({in2[7]} & {in1[5]});
 assign csa_tree_add_55_2_groupi_n_34 = ({in2[1]} & {in1[6]});
 assign csa_tree_add_55_2_groupi_n_33 = ({in2[5]} & {in1[3]});
 assign csa_tree_add_55_2_groupi_n_32 = ({in2[5]} & {in1[5]});
 assign csa_tree_add_55_2_groupi_n_31 = ({in2[0]} & {in1[0]});
 assign csa_tree_add_55_2_groupi_n_30 = ({in2[6]} & {in1[7]});
 assign csa_tree_add_55_2_groupi_n_29 = ({in2[5]} & {in1[7]});
 assign csa_tree_add_55_2_groupi_n_28 = ({in2[0]} & {in1[6]});
 assign csa_tree_add_55_2_groupi_n_27 = ({in2[5]} & {in1[1]});
 assign csa_tree_add_55_2_groupi_n_26 = ({in2[3]} & {in1[1]});
 assign csa_tree_add_55_2_groupi_n_25 = ({in2[1]} & {in1[4]});
 assign csa_tree_add_55_2_groupi_n_24 = ({in2[7]} & {in1[0]});
 assign csa_tree_add_55_2_groupi_n_23 = ({in2[1]} & {in1[0]});
 assign csa_tree_add_55_2_groupi_n_22 = ({in2[4]} & {in1[3]});
 assign csa_tree_add_55_2_groupi_n_21 = ({in2[2]} & {in1[6]});
 assign csa_tree_add_55_2_groupi_n_20 = ({in2[4]} & {in1[6]});
 assign csa_tree_add_55_2_groupi_n_19 = ({in2[3]} & {in1[3]});
 assign csa_tree_add_55_2_groupi_n_18 = ({in2[6]} & {in1[3]});
 assign csa_tree_add_55_2_groupi_n_17 = ({in2[1]} & {in1[2]});
 assign csa_tree_add_55_2_groupi_n_16 = ({in2[6]} & {in1[5]});
 assign csa_tree_add_55_2_groupi_n_15 = ({in2[5]} & {in1[4]});
 assign csa_tree_add_55_2_groupi_n_14 = ({in2[5]} & {in1[0]});
 assign csa_tree_add_55_2_groupi_n_13 = ({in2[1]} & {in1[5]});
 assign csa_tree_add_55_2_groupi_n_12 = ({in2[2]} & {in1[3]});
 assign csa_tree_add_55_2_groupi_n_11 = ({in2[7]} & {in1[4]});
 assign csa_tree_add_55_2_groupi_n_10 = ({in2[4]} & {in1[1]});
 assign csa_tree_add_55_2_groupi_n_9 = ({in2[7]} & {in1[7]});
 assign csa_tree_add_55_2_groupi_n_8 = ({in2[3]} & {in1[6]});
 assign csa_tree_add_55_2_groupi_n_7 = ({in2[3]} & {in1[2]});
 assign csa_tree_add_55_2_groupi_n_6 = ({in2[2]} & {in1[0]});
 assign csa_tree_add_55_2_groupi_n_5 = ({in2[3]} & {in1[4]});
 assign csa_tree_add_55_2_groupi_n_4 = ({in2[4]} & {in1[0]});
 assign csa_tree_add_55_2_groupi_n_3 = ({in2[1]} & {in1[3]});
 assign csa_tree_add_55_2_groupi_n_2 = ({in2[2]} & {in1[7]});
 assign csa_tree_add_55_2_groupi_n_1 = ({in2[7]} & {in1[3]});
 assign csa_tree_add_55_2_groupi_n_0 = ({in2[7]} & {in1[1]});
 assign csa_tree_add_69_2_groupi_n_65 = ~csa_tree_add_69_2_groupi_n_79;
 assign csa_tree_add_69_2_groupi_n_79 = ~n_438;
 assign csa_tree_add_69_2_groupi_n_1583 = ~(csa_tree_add_69_2_groupi_n_1530 & (csa_tree_add_69_2_groupi_n_1582
    | csa_tree_add_69_2_groupi_n_1531));
 assign csa_tree_add_69_2_groupi_n_1582 = ~(csa_tree_add_69_2_groupi_n_1581 | ~csa_tree_add_69_2_groupi_n_1503);
 assign csa_tree_add_69_2_groupi_n_1581 = ~(csa_tree_add_69_2_groupi_n_1567 | csa_tree_add_69_2_groupi_n_1504);
 assign csa_tree_add_69_2_groupi_n_1567 = ~(csa_tree_add_69_2_groupi_n_1557 | csa_tree_add_69_2_groupi_n_58);
 assign csa_tree_add_69_2_groupi_n_1564 = ((csa_tree_add_69_2_groupi_n_1511 & csa_tree_add_69_2_groupi_n_1506)
    | ((csa_tree_add_69_2_groupi_n_1506 & csa_tree_add_69_2_groupi_n_1432) | (csa_tree_add_69_2_groupi_n_1432
    & csa_tree_add_69_2_groupi_n_1511)));
 assign csa_tree_add_69_2_groupi_n_1565 = (csa_tree_add_69_2_groupi_n_1506 ^ (csa_tree_add_69_2_groupi_n_1432
    ^ csa_tree_add_69_2_groupi_n_1511));
 assign csa_tree_add_69_2_groupi_n_1562 = ((csa_tree_add_69_2_groupi_n_1496 & csa_tree_add_69_2_groupi_n_1512)
    | ((csa_tree_add_69_2_groupi_n_1512 & csa_tree_add_69_2_groupi_n_1452) | (csa_tree_add_69_2_groupi_n_1452
    & csa_tree_add_69_2_groupi_n_1496)));
 assign csa_tree_add_69_2_groupi_n_1563 = (csa_tree_add_69_2_groupi_n_1512 ^ (csa_tree_add_69_2_groupi_n_1452
    ^ csa_tree_add_69_2_groupi_n_1496));
 assign csa_tree_add_69_2_groupi_n_1560 = ((csa_tree_add_69_2_groupi_n_1472 & csa_tree_add_69_2_groupi_n_1508)
    | ((csa_tree_add_69_2_groupi_n_1508 & csa_tree_add_69_2_groupi_n_1446) | (csa_tree_add_69_2_groupi_n_1446
    & csa_tree_add_69_2_groupi_n_1472)));
 assign csa_tree_add_69_2_groupi_n_1561 = (csa_tree_add_69_2_groupi_n_1508 ^ (csa_tree_add_69_2_groupi_n_1446
    ^ csa_tree_add_69_2_groupi_n_1472));
 assign csa_tree_add_69_2_groupi_n_1557 = ~(csa_tree_add_69_2_groupi_n_1539 | ~(n_444 | csa_tree_add_69_2_groupi_n_1418));
 assign csa_tree_add_69_2_groupi_n_1555 = ((csa_tree_add_69_2_groupi_n_1507 & csa_tree_add_69_2_groupi_n_1497)
    | ((csa_tree_add_69_2_groupi_n_1497 & csa_tree_add_69_2_groupi_n_1462) | (csa_tree_add_69_2_groupi_n_1462
    & csa_tree_add_69_2_groupi_n_1507)));
 assign csa_tree_add_69_2_groupi_n_1556 = (csa_tree_add_69_2_groupi_n_1497 ^ (csa_tree_add_69_2_groupi_n_1462
    ^ csa_tree_add_69_2_groupi_n_1507));
 assign csa_tree_add_69_2_groupi_n_1548 = ~csa_tree_add_69_2_groupi_n_1539;
 assign csa_tree_add_69_2_groupi_n_1542 = ((csa_tree_add_69_2_groupi_n_1484 & csa_tree_add_69_2_groupi_n_1487)
    | ((csa_tree_add_69_2_groupi_n_1487 & csa_tree_add_69_2_groupi_n_1440) | (csa_tree_add_69_2_groupi_n_1440
    & csa_tree_add_69_2_groupi_n_1484)));
 assign csa_tree_add_69_2_groupi_n_1543 = (csa_tree_add_69_2_groupi_n_1487 ^ (csa_tree_add_69_2_groupi_n_1440
    ^ csa_tree_add_69_2_groupi_n_1484));
 assign csa_tree_add_69_2_groupi_n_1540 = ((csa_tree_add_69_2_groupi_n_1505 & csa_tree_add_69_2_groupi_n_1485)
    | ((csa_tree_add_69_2_groupi_n_1485 & csa_tree_add_69_2_groupi_n_1434) | (csa_tree_add_69_2_groupi_n_1434
    & csa_tree_add_69_2_groupi_n_1505)));
 assign csa_tree_add_69_2_groupi_n_1541 = (csa_tree_add_69_2_groupi_n_1485 ^ (csa_tree_add_69_2_groupi_n_1434
    ^ csa_tree_add_69_2_groupi_n_1505));
 assign csa_tree_add_69_2_groupi_n_1539 = ~(csa_tree_add_69_2_groupi_n_1534 | csa_tree_add_69_2_groupi_n_56);
 assign csa_tree_add_69_2_groupi_n_1537 = ((csa_tree_add_69_2_groupi_n_1473 & csa_tree_add_69_2_groupi_n_1460)
    | ((csa_tree_add_69_2_groupi_n_1460 & csa_tree_add_69_2_groupi_n_1455) | (csa_tree_add_69_2_groupi_n_1455
    & csa_tree_add_69_2_groupi_n_1473)));
 assign csa_tree_add_69_2_groupi_n_1538 = (csa_tree_add_69_2_groupi_n_1460 ^ (csa_tree_add_69_2_groupi_n_1455
    ^ csa_tree_add_69_2_groupi_n_1473));
 assign csa_tree_add_69_2_groupi_n_1535 = ((csa_tree_add_69_2_groupi_n_1429 & csa_tree_add_69_2_groupi_n_1456)
    | ((csa_tree_add_69_2_groupi_n_1456 & csa_tree_add_69_2_groupi_n_1425) | (csa_tree_add_69_2_groupi_n_1425
    & csa_tree_add_69_2_groupi_n_1429)));
 assign csa_tree_add_69_2_groupi_n_1536 = (csa_tree_add_69_2_groupi_n_1456 ^ (csa_tree_add_69_2_groupi_n_1425
    ^ csa_tree_add_69_2_groupi_n_1429));
 assign csa_tree_add_69_2_groupi_n_1534 = ~(csa_tree_add_69_2_groupi_n_1513 | csa_tree_add_69_2_groupi_n_1450);
 assign csa_tree_add_69_2_groupi_n_1533 = ~(csa_tree_add_69_2_groupi_n_1515 ^ csa_tree_add_69_2_groupi_n_1516);
 assign csa_tree_add_69_2_groupi_n_1532 = ~(csa_tree_add_69_2_groupi_n_1529 ^ csa_tree_add_69_2_groupi_n_1500);
 assign csa_tree_add_69_2_groupi_n_1531 = ~(csa_tree_add_69_2_groupi_n_1529 | csa_tree_add_69_2_groupi_n_1500);
 assign csa_tree_add_69_2_groupi_n_1530 = ~(csa_tree_add_69_2_groupi_n_1529 & csa_tree_add_69_2_groupi_n_1500);
 assign csa_tree_add_69_2_groupi_n_1527 = ((csa_tree_add_69_2_groupi_n_1474 & csa_tree_add_69_2_groupi_n_1368)
    | ((csa_tree_add_69_2_groupi_n_1368 & csa_tree_add_69_2_groupi_n_1393) | (csa_tree_add_69_2_groupi_n_1393
    & csa_tree_add_69_2_groupi_n_1474)));
 assign csa_tree_add_69_2_groupi_n_1528 = (csa_tree_add_69_2_groupi_n_1368 ^ (csa_tree_add_69_2_groupi_n_1393
    ^ csa_tree_add_69_2_groupi_n_1474));
 assign csa_tree_add_69_2_groupi_n_1525 = ((csa_tree_add_69_2_groupi_n_1470 & csa_tree_add_69_2_groupi_n_1343)
    | ((csa_tree_add_69_2_groupi_n_1343 & csa_tree_add_69_2_groupi_n_1395) | (csa_tree_add_69_2_groupi_n_1395
    & csa_tree_add_69_2_groupi_n_1470)));
 assign csa_tree_add_69_2_groupi_n_1526 = (csa_tree_add_69_2_groupi_n_1343 ^ (csa_tree_add_69_2_groupi_n_1395
    ^ csa_tree_add_69_2_groupi_n_1470));
 assign csa_tree_add_69_2_groupi_n_1523 = ((csa_tree_add_69_2_groupi_n_1468 & csa_tree_add_69_2_groupi_n_1388)
    | ((csa_tree_add_69_2_groupi_n_1388 & csa_tree_add_69_2_groupi_n_1344) | (csa_tree_add_69_2_groupi_n_1344
    & csa_tree_add_69_2_groupi_n_1468)));
 assign csa_tree_add_69_2_groupi_n_1524 = (csa_tree_add_69_2_groupi_n_1388 ^ (csa_tree_add_69_2_groupi_n_1344
    ^ csa_tree_add_69_2_groupi_n_1468));
 assign csa_tree_add_69_2_groupi_n_1522 = ((csa_tree_add_69_2_groupi_n_1441 & csa_tree_add_69_2_groupi_n_1408)
    | ((csa_tree_add_69_2_groupi_n_1408 & csa_tree_add_69_2_groupi_n_1313) | (csa_tree_add_69_2_groupi_n_1313
    & csa_tree_add_69_2_groupi_n_1441)));
 assign csa_tree_add_69_2_groupi_n_1529 = (csa_tree_add_69_2_groupi_n_1408 ^ (csa_tree_add_69_2_groupi_n_1313
    ^ csa_tree_add_69_2_groupi_n_1441));
 assign csa_tree_add_69_2_groupi_n_1520 = ((csa_tree_add_69_2_groupi_n_1478 & csa_tree_add_69_2_groupi_n_1324)
    | ((csa_tree_add_69_2_groupi_n_1324 & csa_tree_add_69_2_groupi_n_1403) | (csa_tree_add_69_2_groupi_n_1403
    & csa_tree_add_69_2_groupi_n_1478)));
 assign csa_tree_add_69_2_groupi_n_1521 = (csa_tree_add_69_2_groupi_n_1324 ^ (csa_tree_add_69_2_groupi_n_1403
    ^ csa_tree_add_69_2_groupi_n_1478));
 assign csa_tree_add_69_2_groupi_n_1518 = ((csa_tree_add_69_2_groupi_n_1466 & csa_tree_add_69_2_groupi_n_1335)
    | ((csa_tree_add_69_2_groupi_n_1335 & csa_tree_add_69_2_groupi_n_1381) | (csa_tree_add_69_2_groupi_n_1381
    & csa_tree_add_69_2_groupi_n_1466)));
 assign csa_tree_add_69_2_groupi_n_1519 = (csa_tree_add_69_2_groupi_n_1335 ^ (csa_tree_add_69_2_groupi_n_1381
    ^ csa_tree_add_69_2_groupi_n_1466));
 assign csa_tree_add_69_2_groupi_n_1516 = ((csa_tree_add_69_2_groupi_n_1476 & csa_tree_add_69_2_groupi_n_1402)
    | ((csa_tree_add_69_2_groupi_n_1402 & csa_tree_add_69_2_groupi_n_1298) | (csa_tree_add_69_2_groupi_n_1298
    & csa_tree_add_69_2_groupi_n_1476)));
 assign csa_tree_add_69_2_groupi_n_1517 = (csa_tree_add_69_2_groupi_n_1402 ^ (csa_tree_add_69_2_groupi_n_1298
    ^ csa_tree_add_69_2_groupi_n_1476));
 assign csa_tree_add_69_2_groupi_n_1515 = ~(csa_tree_add_69_2_groupi_n_1483 ^ csa_tree_add_69_2_groupi_n_1430);
 assign csa_tree_add_69_2_groupi_n_1514 = ~(csa_tree_add_69_2_groupi_n_1501 ^ csa_tree_add_69_2_groupi_n_1427);
 assign csa_tree_add_69_2_groupi_n_1513 = ~(csa_tree_add_69_2_groupi_n_1502 | csa_tree_add_69_2_groupi_n_53);
 assign csa_tree_add_69_2_groupi_n_1511 = ((csa_tree_add_69_2_groupi_n_1461 & csa_tree_add_69_2_groupi_n_1318)
    | ((csa_tree_add_69_2_groupi_n_1318 & csa_tree_add_69_2_groupi_n_1323) | (csa_tree_add_69_2_groupi_n_1323
    & csa_tree_add_69_2_groupi_n_1461)));
 assign csa_tree_add_69_2_groupi_n_1512 = (csa_tree_add_69_2_groupi_n_1318 ^ (csa_tree_add_69_2_groupi_n_1323
    ^ csa_tree_add_69_2_groupi_n_1461));
 assign csa_tree_add_69_2_groupi_n_1509 = ((csa_tree_add_69_2_groupi_n_1457 & csa_tree_add_69_2_groupi_n_1394)
    | ((csa_tree_add_69_2_groupi_n_1394 & csa_tree_add_69_2_groupi_n_1321) | (csa_tree_add_69_2_groupi_n_1321
    & csa_tree_add_69_2_groupi_n_1457)));
 assign csa_tree_add_69_2_groupi_n_1510 = (csa_tree_add_69_2_groupi_n_1394 ^ (csa_tree_add_69_2_groupi_n_1321
    ^ csa_tree_add_69_2_groupi_n_1457));
 assign csa_tree_add_69_2_groupi_n_1507 = ((csa_tree_add_69_2_groupi_n_1459 & csa_tree_add_69_2_groupi_n_1349)
    | ((csa_tree_add_69_2_groupi_n_1349 & csa_tree_add_69_2_groupi_n_1397) | (csa_tree_add_69_2_groupi_n_1397
    & csa_tree_add_69_2_groupi_n_1459)));
 assign csa_tree_add_69_2_groupi_n_1508 = (csa_tree_add_69_2_groupi_n_1349 ^ (csa_tree_add_69_2_groupi_n_1397
    ^ csa_tree_add_69_2_groupi_n_1459));
 assign csa_tree_add_69_2_groupi_n_1505 = ((csa_tree_add_69_2_groupi_n_1451 & csa_tree_add_69_2_groupi_n_1322)
    | ((csa_tree_add_69_2_groupi_n_1322 & csa_tree_add_69_2_groupi_n_1332) | (csa_tree_add_69_2_groupi_n_1332
    & csa_tree_add_69_2_groupi_n_1451)));
 assign csa_tree_add_69_2_groupi_n_1506 = (csa_tree_add_69_2_groupi_n_1322 ^ (csa_tree_add_69_2_groupi_n_1332
    ^ csa_tree_add_69_2_groupi_n_1451));
 assign csa_tree_add_69_2_groupi_n_1504 = ~(csa_tree_add_69_2_groupi_n_1501 | csa_tree_add_69_2_groupi_n_1427);
 assign csa_tree_add_69_2_groupi_n_1503 = ~(csa_tree_add_69_2_groupi_n_1501 & csa_tree_add_69_2_groupi_n_1427);
 assign csa_tree_add_69_2_groupi_n_1502 = ~(csa_tree_add_69_2_groupi_n_1464 | ~(csa_tree_add_69_2_groupi_n_1407
    | csa_tree_add_69_2_groupi_n_1309));
 assign csa_tree_add_69_2_groupi_n_1498 = ((csa_tree_add_69_2_groupi_n_1447 & csa_tree_add_69_2_groupi_n_1320)
    | ((csa_tree_add_69_2_groupi_n_1320 & csa_tree_add_69_2_groupi_n_1336) | (csa_tree_add_69_2_groupi_n_1336
    & csa_tree_add_69_2_groupi_n_1447)));
 assign csa_tree_add_69_2_groupi_n_1499 = (csa_tree_add_69_2_groupi_n_1320 ^ (csa_tree_add_69_2_groupi_n_1336
    ^ csa_tree_add_69_2_groupi_n_1447));
 assign csa_tree_add_69_2_groupi_n_1496 = ((csa_tree_add_69_2_groupi_n_1445 & csa_tree_add_69_2_groupi_n_1396)
    | ((csa_tree_add_69_2_groupi_n_1396 & csa_tree_add_69_2_groupi_n_1319) | (csa_tree_add_69_2_groupi_n_1319
    & csa_tree_add_69_2_groupi_n_1445)));
 assign csa_tree_add_69_2_groupi_n_1497 = (csa_tree_add_69_2_groupi_n_1396 ^ (csa_tree_add_69_2_groupi_n_1319
    ^ csa_tree_add_69_2_groupi_n_1445));
 assign csa_tree_add_69_2_groupi_n_1494 = ((csa_tree_add_69_2_groupi_n_1443 & csa_tree_add_69_2_groupi_n_1347)
    | ((csa_tree_add_69_2_groupi_n_1347 & csa_tree_add_69_2_groupi_n_1369) | (csa_tree_add_69_2_groupi_n_1369
    & csa_tree_add_69_2_groupi_n_1443)));
 assign csa_tree_add_69_2_groupi_n_1495 = (csa_tree_add_69_2_groupi_n_1347 ^ (csa_tree_add_69_2_groupi_n_1369
    ^ csa_tree_add_69_2_groupi_n_1443));
 assign csa_tree_add_69_2_groupi_n_1500 = ((csa_tree_add_69_2_groupi_n_1442 & csa_tree_add_69_2_groupi_n_1359)
    | ((csa_tree_add_69_2_groupi_n_1359 & csa_tree_add_69_2_groupi_n_1305) | (csa_tree_add_69_2_groupi_n_1305
    & csa_tree_add_69_2_groupi_n_1442)));
 assign csa_tree_add_69_2_groupi_n_1501 = (csa_tree_add_69_2_groupi_n_1359 ^ (csa_tree_add_69_2_groupi_n_1305
    ^ csa_tree_add_69_2_groupi_n_1442));
 assign csa_tree_add_69_2_groupi_n_1492 = ((csa_tree_add_69_2_groupi_n_1435 & csa_tree_add_69_2_groupi_n_1392)
    | ((csa_tree_add_69_2_groupi_n_1392 & csa_tree_add_69_2_groupi_n_1325) | (csa_tree_add_69_2_groupi_n_1325
    & csa_tree_add_69_2_groupi_n_1435)));
 assign csa_tree_add_69_2_groupi_n_1493 = (csa_tree_add_69_2_groupi_n_1392 ^ (csa_tree_add_69_2_groupi_n_1325
    ^ csa_tree_add_69_2_groupi_n_1435));
 assign csa_tree_add_69_2_groupi_n_1490 = ((csa_tree_add_69_2_groupi_n_1439 & csa_tree_add_69_2_groupi_n_1378)
    | ((csa_tree_add_69_2_groupi_n_1378 & csa_tree_add_69_2_groupi_n_1389) | (csa_tree_add_69_2_groupi_n_1389
    & csa_tree_add_69_2_groupi_n_1439)));
 assign csa_tree_add_69_2_groupi_n_1491 = (csa_tree_add_69_2_groupi_n_1378 ^ (csa_tree_add_69_2_groupi_n_1389
    ^ csa_tree_add_69_2_groupi_n_1439));
 assign csa_tree_add_69_2_groupi_n_1488 = ((csa_tree_add_69_2_groupi_n_1437 & csa_tree_add_69_2_groupi_n_1380)
    | ((csa_tree_add_69_2_groupi_n_1380 & csa_tree_add_69_2_groupi_n_1348) | (csa_tree_add_69_2_groupi_n_1348
    & csa_tree_add_69_2_groupi_n_1437)));
 assign csa_tree_add_69_2_groupi_n_1489 = (csa_tree_add_69_2_groupi_n_1380 ^ (csa_tree_add_69_2_groupi_n_1348
    ^ csa_tree_add_69_2_groupi_n_1437));
 assign csa_tree_add_69_2_groupi_n_1486 = ((csa_tree_add_69_2_groupi_n_1433 & csa_tree_add_69_2_groupi_n_1376)
    | ((csa_tree_add_69_2_groupi_n_1376 & csa_tree_add_69_2_groupi_n_1379) | (csa_tree_add_69_2_groupi_n_1379
    & csa_tree_add_69_2_groupi_n_1433)));
 assign csa_tree_add_69_2_groupi_n_1487 = (csa_tree_add_69_2_groupi_n_1376 ^ (csa_tree_add_69_2_groupi_n_1379
    ^ csa_tree_add_69_2_groupi_n_1433));
 assign csa_tree_add_69_2_groupi_n_1484 = ((csa_tree_add_69_2_groupi_n_1431 & csa_tree_add_69_2_groupi_n_1331)
    | ((csa_tree_add_69_2_groupi_n_1331 & csa_tree_add_69_2_groupi_n_1377) | (csa_tree_add_69_2_groupi_n_1377
    & csa_tree_add_69_2_groupi_n_1431)));
 assign csa_tree_add_69_2_groupi_n_1485 = (csa_tree_add_69_2_groupi_n_1331 ^ (csa_tree_add_69_2_groupi_n_1377
    ^ csa_tree_add_69_2_groupi_n_1431));
 assign csa_tree_add_69_2_groupi_n_1483 = ~(csa_tree_add_69_2_groupi_n_1314 ^ csa_tree_add_69_2_groupi_n_1453);
 assign csa_tree_add_69_2_groupi_n_1482 = ~(n_444 ^ csa_tree_add_69_2_groupi_n_1418);
 assign csa_tree_add_69_2_groupi_n_1481 = ~(csa_tree_add_69_2_groupi_n_1413 & (csa_tree_add_69_2_groupi_n_1428
    | csa_tree_add_69_2_groupi_n_1417));
 assign csa_tree_add_69_2_groupi_n_1478 = ((csa_tree_add_69_2_groupi_n_1375 & csa_tree_add_69_2_groupi_n_1111)
    | ((csa_tree_add_69_2_groupi_n_1111 & csa_tree_add_69_2_groupi_n_1386) | (csa_tree_add_69_2_groupi_n_1386
    & csa_tree_add_69_2_groupi_n_1375)));
 assign csa_tree_add_69_2_groupi_n_1479 = (csa_tree_add_69_2_groupi_n_1111 ^ (csa_tree_add_69_2_groupi_n_1386
    ^ csa_tree_add_69_2_groupi_n_1375));
 assign csa_tree_add_69_2_groupi_n_1476 = ((csa_tree_add_69_2_groupi_n_1342 & csa_tree_add_69_2_groupi_n_1148)
    | ((csa_tree_add_69_2_groupi_n_1148 & csa_tree_add_69_2_groupi_n_1374) | (csa_tree_add_69_2_groupi_n_1374
    & csa_tree_add_69_2_groupi_n_1342)));
 assign csa_tree_add_69_2_groupi_n_1477 = (csa_tree_add_69_2_groupi_n_1148 ^ (csa_tree_add_69_2_groupi_n_1374
    ^ csa_tree_add_69_2_groupi_n_1342));
 assign csa_tree_add_69_2_groupi_n_1474 = ((csa_tree_add_69_2_groupi_n_1330 & csa_tree_add_69_2_groupi_n_1123)
    | ((csa_tree_add_69_2_groupi_n_1123 & csa_tree_add_69_2_groupi_n_1398) | (csa_tree_add_69_2_groupi_n_1398
    & csa_tree_add_69_2_groupi_n_1330)));
 assign csa_tree_add_69_2_groupi_n_1475 = (csa_tree_add_69_2_groupi_n_1123 ^ (csa_tree_add_69_2_groupi_n_1398
    ^ csa_tree_add_69_2_groupi_n_1330));
 assign csa_tree_add_69_2_groupi_n_1472 = ((csa_tree_add_69_2_groupi_n_1424 & csa_tree_add_69_2_groupi_n_1306)
    | ((csa_tree_add_69_2_groupi_n_1306 & csa_tree_add_69_2_groupi_n_1350) | (csa_tree_add_69_2_groupi_n_1350
    & csa_tree_add_69_2_groupi_n_1424)));
 assign csa_tree_add_69_2_groupi_n_1473 = (csa_tree_add_69_2_groupi_n_1306 ^ (csa_tree_add_69_2_groupi_n_1350
    ^ csa_tree_add_69_2_groupi_n_1424));
 assign csa_tree_add_69_2_groupi_n_1470 = ((csa_tree_add_69_2_groupi_n_1401 & csa_tree_add_69_2_groupi_n_1129)
    | ((csa_tree_add_69_2_groupi_n_1129 & csa_tree_add_69_2_groupi_n_1384) | (csa_tree_add_69_2_groupi_n_1384
    & csa_tree_add_69_2_groupi_n_1401)));
 assign csa_tree_add_69_2_groupi_n_1471 = (csa_tree_add_69_2_groupi_n_1129 ^ (csa_tree_add_69_2_groupi_n_1384
    ^ csa_tree_add_69_2_groupi_n_1401));
 assign csa_tree_add_69_2_groupi_n_1468 = ((csa_tree_add_69_2_groupi_n_1385 & csa_tree_add_69_2_groupi_n_1179)
    | ((csa_tree_add_69_2_groupi_n_1179 & csa_tree_add_69_2_groupi_n_1382) | (csa_tree_add_69_2_groupi_n_1382
    & csa_tree_add_69_2_groupi_n_1385)));
 assign csa_tree_add_69_2_groupi_n_1469 = (csa_tree_add_69_2_groupi_n_1179 ^ (csa_tree_add_69_2_groupi_n_1382
    ^ csa_tree_add_69_2_groupi_n_1385));
 assign csa_tree_add_69_2_groupi_n_1466 = ((csa_tree_add_69_2_groupi_n_1338 & csa_tree_add_69_2_groupi_n_1113)
    | ((csa_tree_add_69_2_groupi_n_1113 & csa_tree_add_69_2_groupi_n_1372) | (csa_tree_add_69_2_groupi_n_1372
    & csa_tree_add_69_2_groupi_n_1338)));
 assign csa_tree_add_69_2_groupi_n_1467 = (csa_tree_add_69_2_groupi_n_1113 ^ (csa_tree_add_69_2_groupi_n_1372
    ^ csa_tree_add_69_2_groupi_n_1338));
 assign csa_tree_add_69_2_groupi_n_1463 = ~(n_445 ^ csa_tree_add_69_2_groupi_n_1406);
 assign csa_tree_add_69_2_groupi_n_1464 = ~(csa_tree_add_69_2_groupi_n_1449 | csa_tree_add_69_2_groupi_n_51);
 assign csa_tree_add_69_2_groupi_n_1461 = ((csa_tree_add_69_2_groupi_n_1367 & csa_tree_add_69_2_groupi_n_1165)
    | ((csa_tree_add_69_2_groupi_n_1165 & csa_tree_add_69_2_groupi_n_1355) | (csa_tree_add_69_2_groupi_n_1355
    & csa_tree_add_69_2_groupi_n_1367)));
 assign csa_tree_add_69_2_groupi_n_1462 = (csa_tree_add_69_2_groupi_n_1165 ^ (csa_tree_add_69_2_groupi_n_1355
    ^ csa_tree_add_69_2_groupi_n_1367));
 assign csa_tree_add_69_2_groupi_n_1459 = ((csa_tree_add_69_2_groupi_n_1390 & csa_tree_add_69_2_groupi_n_1175)
    | ((csa_tree_add_69_2_groupi_n_1175 & csa_tree_add_69_2_groupi_n_1352) | (csa_tree_add_69_2_groupi_n_1352
    & csa_tree_add_69_2_groupi_n_1390)));
 assign csa_tree_add_69_2_groupi_n_1460 = (csa_tree_add_69_2_groupi_n_1175 ^ (csa_tree_add_69_2_groupi_n_1352
    ^ csa_tree_add_69_2_groupi_n_1390));
 assign csa_tree_add_69_2_groupi_n_1457 = ((csa_tree_add_69_2_groupi_n_1400 & csa_tree_add_69_2_groupi_n_1117)
    | ((csa_tree_add_69_2_groupi_n_1117 & csa_tree_add_69_2_groupi_n_1354) | (csa_tree_add_69_2_groupi_n_1354
    & csa_tree_add_69_2_groupi_n_1400)));
 assign csa_tree_add_69_2_groupi_n_1458 = (csa_tree_add_69_2_groupi_n_1117 ^ (csa_tree_add_69_2_groupi_n_1354
    ^ csa_tree_add_69_2_groupi_n_1400));
 assign csa_tree_add_69_2_groupi_n_1455 = ((csa_tree_add_69_2_groupi_n_1410 & csa_tree_add_69_2_groupi_n_1283)
    | ((csa_tree_add_69_2_groupi_n_1283 & csa_tree_add_69_2_groupi_n_1307) | (csa_tree_add_69_2_groupi_n_1307
    & csa_tree_add_69_2_groupi_n_1410)));
 assign csa_tree_add_69_2_groupi_n_1456 = (csa_tree_add_69_2_groupi_n_1283 ^ (csa_tree_add_69_2_groupi_n_1307
    ^ csa_tree_add_69_2_groupi_n_1410));
 assign csa_tree_add_69_2_groupi_n_1453 = ((csa_tree_add_69_2_groupi_n_1371 & csa_tree_add_69_2_groupi_n_1150)
    | ((csa_tree_add_69_2_groupi_n_1150 & csa_tree_add_69_2_groupi_n_1341) | (csa_tree_add_69_2_groupi_n_1341
    & csa_tree_add_69_2_groupi_n_1371)));
 assign csa_tree_add_69_2_groupi_n_1454 = (csa_tree_add_69_2_groupi_n_1150 ^ (csa_tree_add_69_2_groupi_n_1341
    ^ csa_tree_add_69_2_groupi_n_1371));
 assign csa_tree_add_69_2_groupi_n_1451 = ((csa_tree_add_69_2_groupi_n_1366 & csa_tree_add_69_2_groupi_n_1125)
    | ((csa_tree_add_69_2_groupi_n_1125 & csa_tree_add_69_2_groupi_n_1328) | (csa_tree_add_69_2_groupi_n_1328
    & csa_tree_add_69_2_groupi_n_1366)));
 assign csa_tree_add_69_2_groupi_n_1452 = (csa_tree_add_69_2_groupi_n_1125 ^ (csa_tree_add_69_2_groupi_n_1328
    ^ csa_tree_add_69_2_groupi_n_1366));
 assign csa_tree_add_69_2_groupi_n_1450 = ~(n_445 | csa_tree_add_69_2_groupi_n_1406);
 assign csa_tree_add_69_2_groupi_n_1449 = ~(csa_tree_add_69_2_groupi_n_1420 | ~(n_446 | csa_tree_add_69_2_groupi_n_1310));
 assign csa_tree_add_69_2_groupi_n_1447 = ((csa_tree_add_69_2_groupi_n_1353 & csa_tree_add_69_2_groupi_n_1115)
    | ((csa_tree_add_69_2_groupi_n_1115 & csa_tree_add_69_2_groupi_n_1373) | (csa_tree_add_69_2_groupi_n_1373
    & csa_tree_add_69_2_groupi_n_1353)));
 assign csa_tree_add_69_2_groupi_n_1448 = (csa_tree_add_69_2_groupi_n_1115 ^ (csa_tree_add_69_2_groupi_n_1373
    ^ csa_tree_add_69_2_groupi_n_1353));
 assign csa_tree_add_69_2_groupi_n_1445 = ((csa_tree_add_69_2_groupi_n_1351 & csa_tree_add_69_2_groupi_n_1121)
    | ((csa_tree_add_69_2_groupi_n_1121 & csa_tree_add_69_2_groupi_n_1356) | (csa_tree_add_69_2_groupi_n_1356
    & csa_tree_add_69_2_groupi_n_1351)));
 assign csa_tree_add_69_2_groupi_n_1446 = (csa_tree_add_69_2_groupi_n_1121 ^ (csa_tree_add_69_2_groupi_n_1356
    ^ csa_tree_add_69_2_groupi_n_1351));
 assign csa_tree_add_69_2_groupi_n_1443 = ((csa_tree_add_69_2_groupi_n_1339 & csa_tree_add_69_2_groupi_n_1156)
    | ((csa_tree_add_69_2_groupi_n_1156 & csa_tree_add_69_2_groupi_n_1399) | (csa_tree_add_69_2_groupi_n_1399
    & csa_tree_add_69_2_groupi_n_1339)));
 assign csa_tree_add_69_2_groupi_n_1444 = (csa_tree_add_69_2_groupi_n_1156 ^ (csa_tree_add_69_2_groupi_n_1399
    ^ csa_tree_add_69_2_groupi_n_1339));
 assign csa_tree_add_69_2_groupi_n_1441 = ((csa_tree_add_69_2_groupi_n_1326 & csa_tree_add_69_2_groupi_n_1284)
    | ((csa_tree_add_69_2_groupi_n_1284 & csa_tree_add_69_2_groupi_n_1089) | (csa_tree_add_69_2_groupi_n_1089
    & csa_tree_add_69_2_groupi_n_1326)));
 assign csa_tree_add_69_2_groupi_n_1442 = (csa_tree_add_69_2_groupi_n_1284 ^ (csa_tree_add_69_2_groupi_n_1089
    ^ csa_tree_add_69_2_groupi_n_1326));
 assign csa_tree_add_69_2_groupi_n_1439 = ((csa_tree_add_69_2_groupi_n_1345 & csa_tree_add_69_2_groupi_n_1187)
    | ((csa_tree_add_69_2_groupi_n_1187 & csa_tree_add_69_2_groupi_n_1383) | (csa_tree_add_69_2_groupi_n_1383
    & csa_tree_add_69_2_groupi_n_1345)));
 assign csa_tree_add_69_2_groupi_n_1440 = (csa_tree_add_69_2_groupi_n_1187 ^ (csa_tree_add_69_2_groupi_n_1383
    ^ csa_tree_add_69_2_groupi_n_1345));
 assign csa_tree_add_69_2_groupi_n_1437 = ((csa_tree_add_69_2_groupi_n_1337 & csa_tree_add_69_2_groupi_n_1127)
    | ((csa_tree_add_69_2_groupi_n_1127 & csa_tree_add_69_2_groupi_n_1340) | (csa_tree_add_69_2_groupi_n_1340
    & csa_tree_add_69_2_groupi_n_1337)));
 assign csa_tree_add_69_2_groupi_n_1438 = (csa_tree_add_69_2_groupi_n_1127 ^ (csa_tree_add_69_2_groupi_n_1340
    ^ csa_tree_add_69_2_groupi_n_1337));
 assign csa_tree_add_69_2_groupi_n_1435 = ((csa_tree_add_69_2_groupi_n_1329 & csa_tree_add_69_2_groupi_n_1135)
    | ((csa_tree_add_69_2_groupi_n_1135 & csa_tree_add_69_2_groupi_n_1387) | (csa_tree_add_69_2_groupi_n_1387
    & csa_tree_add_69_2_groupi_n_1329)));
 assign csa_tree_add_69_2_groupi_n_1436 = (csa_tree_add_69_2_groupi_n_1135 ^ (csa_tree_add_69_2_groupi_n_1387
    ^ csa_tree_add_69_2_groupi_n_1329));
 assign csa_tree_add_69_2_groupi_n_1433 = ((csa_tree_add_69_2_groupi_n_1333 & csa_tree_add_69_2_groupi_n_1109)
    | ((csa_tree_add_69_2_groupi_n_1109 & csa_tree_add_69_2_groupi_n_1346) | (csa_tree_add_69_2_groupi_n_1346
    & csa_tree_add_69_2_groupi_n_1333)));
 assign csa_tree_add_69_2_groupi_n_1434 = (csa_tree_add_69_2_groupi_n_1109 ^ (csa_tree_add_69_2_groupi_n_1346
    ^ csa_tree_add_69_2_groupi_n_1333));
 assign csa_tree_add_69_2_groupi_n_1431 = ((csa_tree_add_69_2_groupi_n_1327 & csa_tree_add_69_2_groupi_n_1173)
    | ((csa_tree_add_69_2_groupi_n_1173 & csa_tree_add_69_2_groupi_n_1334) | (csa_tree_add_69_2_groupi_n_1334
    & csa_tree_add_69_2_groupi_n_1327)));
 assign csa_tree_add_69_2_groupi_n_1432 = (csa_tree_add_69_2_groupi_n_1173 ^ (csa_tree_add_69_2_groupi_n_1334
    ^ csa_tree_add_69_2_groupi_n_1327));
 assign csa_tree_add_69_2_groupi_n_1430 = ~(csa_tree_add_69_2_groupi_n_1412 ^ csa_tree_add_69_2_groupi_n_1290);
 assign csa_tree_add_69_2_groupi_n_1429 = ~(csa_tree_add_69_2_groupi_n_1365 & (csa_tree_add_69_2_groupi_n_1363
    | csa_tree_add_69_2_groupi_n_1315));
 assign csa_tree_add_69_2_groupi_n_1428 = ~(csa_tree_add_69_2_groupi_n_1404 ^ csa_tree_add_69_2_groupi_n_1315);
 assign csa_tree_add_69_2_groupi_n_1427 = ~(csa_tree_add_69_2_groupi_n_1362 & (csa_tree_add_69_2_groupi_n_93
    | csa_tree_add_69_2_groupi_n_1364));
 assign csa_tree_add_69_2_groupi_n_1424 = ((csa_tree_add_69_2_groupi_n_1391 & csa_tree_add_69_2_groupi_n_1191)
    | ((csa_tree_add_69_2_groupi_n_1191 & csa_tree_add_69_2_groupi_n_1299) | (csa_tree_add_69_2_groupi_n_1299
    & csa_tree_add_69_2_groupi_n_1391)));
 assign csa_tree_add_69_2_groupi_n_1425 = (csa_tree_add_69_2_groupi_n_1191 ^ (csa_tree_add_69_2_groupi_n_1299
    ^ csa_tree_add_69_2_groupi_n_1391));
 assign csa_tree_add_69_2_groupi_n_1421 = ~(csa_tree_add_69_2_groupi_n_1407 ^ csa_tree_add_69_2_groupi_n_1309);
 assign csa_tree_add_69_2_groupi_n_1420 = ~(csa_tree_add_69_2_groupi_n_1414 | csa_tree_add_69_2_groupi_n_50);
 assign csa_tree_add_69_2_groupi_n_1418 = ~(csa_tree_add_69_2_groupi_n_1316 & (csa_tree_add_69_2_groupi_n_1303
    | csa_tree_add_69_2_groupi_n_1317));
 assign csa_tree_add_69_2_groupi_n_1417 = ~(csa_tree_add_69_2_groupi_n_1411 | csa_tree_add_69_2_groupi_n_1409);
 assign csa_tree_add_69_2_groupi_n_1414 = ~(csa_tree_add_69_2_groupi_n_1294 | ~(csa_tree_add_69_2_groupi_n_1311
    | csa_tree_add_69_2_groupi_n_1214));
 assign csa_tree_add_69_2_groupi_n_1413 = ~(csa_tree_add_69_2_groupi_n_1411 & csa_tree_add_69_2_groupi_n_1409);
 assign csa_tree_add_69_2_groupi_n_1412 = ~(csa_tree_add_69_2_groupi_n_1077 ^ csa_tree_add_69_2_groupi_n_1370);
 assign csa_tree_add_69_2_groupi_n_1410 = ((csa_tree_add_69_2_groupi_n_1300 & csa_tree_add_69_2_groupi_n_1105)
    | ((csa_tree_add_69_2_groupi_n_1105 & csa_tree_add_69_2_groupi_n_1270) | (csa_tree_add_69_2_groupi_n_1270
    & csa_tree_add_69_2_groupi_n_1300)));
 assign csa_tree_add_69_2_groupi_n_1411 = (csa_tree_add_69_2_groupi_n_1105 ^ (csa_tree_add_69_2_groupi_n_1270
    ^ csa_tree_add_69_2_groupi_n_1300));
 assign csa_tree_add_69_2_groupi_n_1409 = ((csa_tree_add_69_2_groupi_n_1304 & csa_tree_add_69_2_groupi_n_44)
    | ((csa_tree_add_69_2_groupi_n_44 & csa_tree_add_69_2_groupi_n_1271) | (csa_tree_add_69_2_groupi_n_1271
    & csa_tree_add_69_2_groupi_n_1304)));
 assign csa_tree_add_69_2_groupi_n_1408 = (csa_tree_add_69_2_groupi_n_44 ^ (csa_tree_add_69_2_groupi_n_1271
    ^ csa_tree_add_69_2_groupi_n_1304));
 assign csa_tree_add_69_2_groupi_n_1406 = ((csa_tree_add_69_2_groupi_n_1293 & csa_tree_add_69_2_groupi_n_1215)
    | ((csa_tree_add_69_2_groupi_n_1215 & csa_tree_add_69_2_groupi_n_1075) | (csa_tree_add_69_2_groupi_n_1075
    & csa_tree_add_69_2_groupi_n_1293)));
 assign csa_tree_add_69_2_groupi_n_1407 = (csa_tree_add_69_2_groupi_n_1215 ^ (csa_tree_add_69_2_groupi_n_1075
    ^ csa_tree_add_69_2_groupi_n_1293));
 assign csa_tree_add_69_2_groupi_n_1405 = ~(n_446 ^ csa_tree_add_69_2_groupi_n_1310);
 assign csa_tree_add_69_2_groupi_n_1404 = ~((csa_tree_add_69_2_groupi_n_1218 & ~csa_tree_add_69_2_groupi_n_1308)
    | (csa_tree_add_69_2_groupi_n_1280 & csa_tree_add_69_2_groupi_n_1308));
 assign csa_tree_add_69_2_groupi_n_1402 = ((csa_tree_add_69_2_groupi_n_1262 & csa_tree_add_69_2_groupi_n_1110)
    | ((csa_tree_add_69_2_groupi_n_1110 & csa_tree_add_69_2_groupi_n_1162) | (csa_tree_add_69_2_groupi_n_1162
    & csa_tree_add_69_2_groupi_n_1262)));
 assign csa_tree_add_69_2_groupi_n_1403 = (csa_tree_add_69_2_groupi_n_1110 ^ (csa_tree_add_69_2_groupi_n_1162
    ^ csa_tree_add_69_2_groupi_n_1262));
 assign csa_tree_add_69_2_groupi_n_1400 = ((csa_tree_add_69_2_groupi_n_1276 & csa_tree_add_69_2_groupi_n_1159)
    | ((csa_tree_add_69_2_groupi_n_1159 & csa_tree_add_69_2_groupi_n_895) | (csa_tree_add_69_2_groupi_n_895
    & csa_tree_add_69_2_groupi_n_1276)));
 assign csa_tree_add_69_2_groupi_n_1401 = (csa_tree_add_69_2_groupi_n_1159 ^ (csa_tree_add_69_2_groupi_n_895
    ^ csa_tree_add_69_2_groupi_n_1276));
 assign csa_tree_add_69_2_groupi_n_1398 = ((csa_tree_add_69_2_groupi_n_1259 & csa_tree_add_69_2_groupi_n_1098)
    | ((csa_tree_add_69_2_groupi_n_1098 & csa_tree_add_69_2_groupi_n_892) | (csa_tree_add_69_2_groupi_n_892
    & csa_tree_add_69_2_groupi_n_1259)));
 assign csa_tree_add_69_2_groupi_n_1399 = (csa_tree_add_69_2_groupi_n_1098 ^ (csa_tree_add_69_2_groupi_n_892
    ^ csa_tree_add_69_2_groupi_n_1259));
 assign csa_tree_add_69_2_groupi_n_1396 = ((csa_tree_add_69_2_groupi_n_1264 & csa_tree_add_69_2_groupi_n_1174)
    | ((csa_tree_add_69_2_groupi_n_1174 & csa_tree_add_69_2_groupi_n_1181) | (csa_tree_add_69_2_groupi_n_1181
    & csa_tree_add_69_2_groupi_n_1264)));
 assign csa_tree_add_69_2_groupi_n_1397 = (csa_tree_add_69_2_groupi_n_1174 ^ (csa_tree_add_69_2_groupi_n_1181
    ^ csa_tree_add_69_2_groupi_n_1264));
 assign csa_tree_add_69_2_groupi_n_1394 = ((csa_tree_add_69_2_groupi_n_1266 & csa_tree_add_69_2_groupi_n_1128)
    | ((csa_tree_add_69_2_groupi_n_1128 & csa_tree_add_69_2_groupi_n_1131) | (csa_tree_add_69_2_groupi_n_1131
    & csa_tree_add_69_2_groupi_n_1266)));
 assign csa_tree_add_69_2_groupi_n_1395 = (csa_tree_add_69_2_groupi_n_1128 ^ (csa_tree_add_69_2_groupi_n_1131
    ^ csa_tree_add_69_2_groupi_n_1266));
 assign csa_tree_add_69_2_groupi_n_1392 = ((csa_tree_add_69_2_groupi_n_1275 & csa_tree_add_69_2_groupi_n_1122)
    | ((csa_tree_add_69_2_groupi_n_1122 & csa_tree_add_69_2_groupi_n_1189) | (csa_tree_add_69_2_groupi_n_1189
    & csa_tree_add_69_2_groupi_n_1275)));
 assign csa_tree_add_69_2_groupi_n_1393 = (csa_tree_add_69_2_groupi_n_1122 ^ (csa_tree_add_69_2_groupi_n_1189
    ^ csa_tree_add_69_2_groupi_n_1275));
 assign csa_tree_add_69_2_groupi_n_1390 = ((csa_tree_add_69_2_groupi_n_1245 & csa_tree_add_69_2_groupi_n_900)
    | ((csa_tree_add_69_2_groupi_n_900 & csa_tree_add_69_2_groupi_n_1242) | (csa_tree_add_69_2_groupi_n_1242
    & csa_tree_add_69_2_groupi_n_1245)));
 assign csa_tree_add_69_2_groupi_n_1391 = (csa_tree_add_69_2_groupi_n_900 ^ (csa_tree_add_69_2_groupi_n_1242
    ^ csa_tree_add_69_2_groupi_n_1245));
 assign csa_tree_add_69_2_groupi_n_1388 = ((csa_tree_add_69_2_groupi_n_1277 & csa_tree_add_69_2_groupi_n_1186)
    | ((csa_tree_add_69_2_groupi_n_1186 & csa_tree_add_69_2_groupi_n_1160) | (csa_tree_add_69_2_groupi_n_1160
    & csa_tree_add_69_2_groupi_n_1277)));
 assign csa_tree_add_69_2_groupi_n_1389 = (csa_tree_add_69_2_groupi_n_1186 ^ (csa_tree_add_69_2_groupi_n_1160
    ^ csa_tree_add_69_2_groupi_n_1277));
 assign csa_tree_add_69_2_groupi_n_1386 = ((csa_tree_add_69_2_groupi_n_1278 & csa_tree_add_69_2_groupi_n_1166)
    | ((csa_tree_add_69_2_groupi_n_1166 & csa_tree_add_69_2_groupi_n_918) | (csa_tree_add_69_2_groupi_n_918
    & csa_tree_add_69_2_groupi_n_1278)));
 assign csa_tree_add_69_2_groupi_n_1387 = (csa_tree_add_69_2_groupi_n_1166 ^ (csa_tree_add_69_2_groupi_n_918
    ^ csa_tree_add_69_2_groupi_n_1278));
 assign csa_tree_add_69_2_groupi_n_1384 = ((csa_tree_add_69_2_groupi_n_1272 & csa_tree_add_69_2_groupi_n_1182)
    | ((csa_tree_add_69_2_groupi_n_1182 & csa_tree_add_69_2_groupi_n_917) | (csa_tree_add_69_2_groupi_n_917
    & csa_tree_add_69_2_groupi_n_1272)));
 assign csa_tree_add_69_2_groupi_n_1385 = (csa_tree_add_69_2_groupi_n_1182 ^ (csa_tree_add_69_2_groupi_n_917
    ^ csa_tree_add_69_2_groupi_n_1272));
 assign csa_tree_add_69_2_groupi_n_1382 = ((csa_tree_add_69_2_groupi_n_1267 & csa_tree_add_69_2_groupi_n_1151)
    | ((csa_tree_add_69_2_groupi_n_1151 & csa_tree_add_69_2_groupi_n_882) | (csa_tree_add_69_2_groupi_n_882
    & csa_tree_add_69_2_groupi_n_1267)));
 assign csa_tree_add_69_2_groupi_n_1383 = (csa_tree_add_69_2_groupi_n_1151 ^ (csa_tree_add_69_2_groupi_n_882
    ^ csa_tree_add_69_2_groupi_n_1267));
 assign csa_tree_add_69_2_groupi_n_1380 = ((csa_tree_add_69_2_groupi_n_1260 & csa_tree_add_69_2_groupi_n_1112)
    | ((csa_tree_add_69_2_groupi_n_1112 & csa_tree_add_69_2_groupi_n_1099) | (csa_tree_add_69_2_groupi_n_1099
    & csa_tree_add_69_2_groupi_n_1260)));
 assign csa_tree_add_69_2_groupi_n_1381 = (csa_tree_add_69_2_groupi_n_1112 ^ (csa_tree_add_69_2_groupi_n_1099
    ^ csa_tree_add_69_2_groupi_n_1260));
 assign csa_tree_add_69_2_groupi_n_1378 = ((csa_tree_add_69_2_groupi_n_1273 & csa_tree_add_69_2_groupi_n_1108)
    | ((csa_tree_add_69_2_groupi_n_1108 & csa_tree_add_69_2_groupi_n_1183) | (csa_tree_add_69_2_groupi_n_1183
    & csa_tree_add_69_2_groupi_n_1273)));
 assign csa_tree_add_69_2_groupi_n_1379 = (csa_tree_add_69_2_groupi_n_1108 ^ (csa_tree_add_69_2_groupi_n_1183
    ^ csa_tree_add_69_2_groupi_n_1273));
 assign csa_tree_add_69_2_groupi_n_1376 = ((csa_tree_add_69_2_groupi_n_1268 & csa_tree_add_69_2_groupi_n_1172)
    | ((csa_tree_add_69_2_groupi_n_1172 & csa_tree_add_69_2_groupi_n_1152) | (csa_tree_add_69_2_groupi_n_1152
    & csa_tree_add_69_2_groupi_n_1268)));
 assign csa_tree_add_69_2_groupi_n_1377 = (csa_tree_add_69_2_groupi_n_1172 ^ (csa_tree_add_69_2_groupi_n_1152
    ^ csa_tree_add_69_2_groupi_n_1268));
 assign csa_tree_add_69_2_groupi_n_1374 = ((csa_tree_add_69_2_groupi_n_1274 & csa_tree_add_69_2_groupi_n_1188)
    | ((csa_tree_add_69_2_groupi_n_1188 & csa_tree_add_69_2_groupi_n_894) | (csa_tree_add_69_2_groupi_n_894
    & csa_tree_add_69_2_groupi_n_1274)));
 assign csa_tree_add_69_2_groupi_n_1375 = (csa_tree_add_69_2_groupi_n_1188 ^ (csa_tree_add_69_2_groupi_n_894
    ^ csa_tree_add_69_2_groupi_n_1274));
 assign csa_tree_add_69_2_groupi_n_1372 = ((csa_tree_add_69_2_groupi_n_1265 & csa_tree_add_69_2_groupi_n_1130)
    | ((csa_tree_add_69_2_groupi_n_1130 & csa_tree_add_69_2_groupi_n_912) | (csa_tree_add_69_2_groupi_n_912
    & csa_tree_add_69_2_groupi_n_1265)));
 assign csa_tree_add_69_2_groupi_n_1373 = (csa_tree_add_69_2_groupi_n_1130 ^ (csa_tree_add_69_2_groupi_n_912
    ^ csa_tree_add_69_2_groupi_n_1265));
 assign csa_tree_add_69_2_groupi_n_1370 = ((csa_tree_add_69_2_groupi_n_1261 & csa_tree_add_69_2_groupi_n_1154)
    | ((csa_tree_add_69_2_groupi_n_1154 & csa_tree_add_69_2_groupi_n_887) | (csa_tree_add_69_2_groupi_n_887
    & csa_tree_add_69_2_groupi_n_1261)));
 assign csa_tree_add_69_2_groupi_n_1371 = (csa_tree_add_69_2_groupi_n_1154 ^ (csa_tree_add_69_2_groupi_n_887
    ^ csa_tree_add_69_2_groupi_n_1261));
 assign csa_tree_add_69_2_groupi_n_1368 = ((csa_tree_add_69_2_groupi_n_1279 & csa_tree_add_69_2_groupi_n_1155)
    | ((csa_tree_add_69_2_groupi_n_1155 & csa_tree_add_69_2_groupi_n_1167) | (csa_tree_add_69_2_groupi_n_1167
    & csa_tree_add_69_2_groupi_n_1279)));
 assign csa_tree_add_69_2_groupi_n_1369 = (csa_tree_add_69_2_groupi_n_1155 ^ (csa_tree_add_69_2_groupi_n_1167
    ^ csa_tree_add_69_2_groupi_n_1279));
 assign csa_tree_add_69_2_groupi_n_1366 = ((csa_tree_add_69_2_groupi_n_1263 & csa_tree_add_69_2_groupi_n_1180)
    | ((csa_tree_add_69_2_groupi_n_1180 & csa_tree_add_69_2_groupi_n_914) | (csa_tree_add_69_2_groupi_n_914
    & csa_tree_add_69_2_groupi_n_1263)));
 assign csa_tree_add_69_2_groupi_n_1367 = (csa_tree_add_69_2_groupi_n_1180 ^ (csa_tree_add_69_2_groupi_n_914
    ^ csa_tree_add_69_2_groupi_n_1263));
 assign csa_tree_add_69_2_groupi_n_1365 = ~(csa_tree_add_69_2_groupi_n_1358 & csa_tree_add_69_2_groupi_n_1280);
 assign csa_tree_add_69_2_groupi_n_1364 = ~(csa_tree_add_69_2_groupi_n_1357 | csa_tree_add_69_2_groupi_n_1287);
 assign csa_tree_add_69_2_groupi_n_1363 = ~(csa_tree_add_69_2_groupi_n_1358 | csa_tree_add_69_2_groupi_n_1280);
 assign csa_tree_add_69_2_groupi_n_1362 = ~(csa_tree_add_69_2_groupi_n_1357 & csa_tree_add_69_2_groupi_n_1287);
 assign csa_tree_add_69_2_groupi_n_1360 = ~(csa_tree_add_69_2_groupi_n_1311 ^ csa_tree_add_69_2_groupi_n_1214);
 assign csa_tree_add_69_2_groupi_n_1361 = ~((csa_tree_add_69_2_groupi_n_1301 & ~csa_tree_add_69_2_groupi_n_1286)
    | (csa_tree_add_69_2_groupi_n_1312 & csa_tree_add_69_2_groupi_n_1286));
 assign csa_tree_add_69_2_groupi_n_1359 = ~((csa_tree_add_69_2_groupi_n_1288 & csa_tree_add_69_2_groupi_n_1282)
    | ((csa_tree_add_69_2_groupi_n_1282 & csa_tree_add_69_2_groupi_n_1201) | (csa_tree_add_69_2_groupi_n_1201
    & csa_tree_add_69_2_groupi_n_1288)));
 assign csa_tree_add_69_2_groupi_n_1358 = ~csa_tree_add_69_2_groupi_n_1308;
 assign csa_tree_add_69_2_groupi_n_1355 = ((csa_tree_add_69_2_groupi_n_1225 & csa_tree_add_69_2_groupi_n_1170)
    | ((csa_tree_add_69_2_groupi_n_1170 & csa_tree_add_69_2_groupi_n_910) | (csa_tree_add_69_2_groupi_n_910
    & csa_tree_add_69_2_groupi_n_1225)));
 assign csa_tree_add_69_2_groupi_n_1356 = (csa_tree_add_69_2_groupi_n_1170 ^ (csa_tree_add_69_2_groupi_n_910
    ^ csa_tree_add_69_2_groupi_n_1225));
 assign csa_tree_add_69_2_groupi_n_1353 = ((csa_tree_add_69_2_groupi_n_1227 & csa_tree_add_69_2_groupi_n_1145)
    | ((csa_tree_add_69_2_groupi_n_1145 & csa_tree_add_69_2_groupi_n_902) | (csa_tree_add_69_2_groupi_n_902
    & csa_tree_add_69_2_groupi_n_1227)));
 assign csa_tree_add_69_2_groupi_n_1354 = (csa_tree_add_69_2_groupi_n_1145 ^ (csa_tree_add_69_2_groupi_n_902
    ^ csa_tree_add_69_2_groupi_n_1227));
 assign csa_tree_add_69_2_groupi_n_1351 = ((csa_tree_add_69_2_groupi_n_1244 & csa_tree_add_69_2_groupi_n_1132)
    | ((csa_tree_add_69_2_groupi_n_1132 & csa_tree_add_69_2_groupi_n_905) | (csa_tree_add_69_2_groupi_n_905
    & csa_tree_add_69_2_groupi_n_1244)));
 assign csa_tree_add_69_2_groupi_n_1352 = (csa_tree_add_69_2_groupi_n_1132 ^ (csa_tree_add_69_2_groupi_n_905
    ^ csa_tree_add_69_2_groupi_n_1244));
 assign csa_tree_add_69_2_groupi_n_1349 = ((csa_tree_add_69_2_groupi_n_1226 & csa_tree_add_69_2_groupi_n_1190)
    | ((csa_tree_add_69_2_groupi_n_1190 & csa_tree_add_69_2_groupi_n_1171) | (csa_tree_add_69_2_groupi_n_1171
    & csa_tree_add_69_2_groupi_n_1226)));
 assign csa_tree_add_69_2_groupi_n_1350 = (csa_tree_add_69_2_groupi_n_1190 ^ (csa_tree_add_69_2_groupi_n_1171
    ^ csa_tree_add_69_2_groupi_n_1226));
 assign csa_tree_add_69_2_groupi_n_1347 = ((csa_tree_add_69_2_groupi_n_1239 & csa_tree_add_69_2_groupi_n_1126)
    | ((csa_tree_add_69_2_groupi_n_1126 & csa_tree_add_69_2_groupi_n_1103) | (csa_tree_add_69_2_groupi_n_1103
    & csa_tree_add_69_2_groupi_n_1239)));
 assign csa_tree_add_69_2_groupi_n_1348 = (csa_tree_add_69_2_groupi_n_1126 ^ (csa_tree_add_69_2_groupi_n_1103
    ^ csa_tree_add_69_2_groupi_n_1239));
 assign csa_tree_add_69_2_groupi_n_1345 = ((csa_tree_add_69_2_groupi_n_1246 & csa_tree_add_69_2_groupi_n_1157)
    | ((csa_tree_add_69_2_groupi_n_1157 & csa_tree_add_69_2_groupi_n_883) | (csa_tree_add_69_2_groupi_n_883
    & csa_tree_add_69_2_groupi_n_1246)));
 assign csa_tree_add_69_2_groupi_n_1346 = (csa_tree_add_69_2_groupi_n_1157 ^ (csa_tree_add_69_2_groupi_n_883
    ^ csa_tree_add_69_2_groupi_n_1246));
 assign csa_tree_add_69_2_groupi_n_1343 = ((csa_tree_add_69_2_groupi_n_1228 & csa_tree_add_69_2_groupi_n_1178)
    | ((csa_tree_add_69_2_groupi_n_1178 & csa_tree_add_69_2_groupi_n_1146) | (csa_tree_add_69_2_groupi_n_1146
    & csa_tree_add_69_2_groupi_n_1228)));
 assign csa_tree_add_69_2_groupi_n_1344 = (csa_tree_add_69_2_groupi_n_1178 ^ (csa_tree_add_69_2_groupi_n_1146
    ^ csa_tree_add_69_2_groupi_n_1228));
 assign csa_tree_add_69_2_groupi_n_1341 = ((csa_tree_add_69_2_groupi_n_1234 & csa_tree_add_69_2_groupi_n_1184)
    | ((csa_tree_add_69_2_groupi_n_1184 & csa_tree_add_69_2_groupi_n_888) | (csa_tree_add_69_2_groupi_n_888
    & csa_tree_add_69_2_groupi_n_1234)));
 assign csa_tree_add_69_2_groupi_n_1342 = (csa_tree_add_69_2_groupi_n_1184 ^ (csa_tree_add_69_2_groupi_n_888
    ^ csa_tree_add_69_2_groupi_n_1234));
 assign csa_tree_add_69_2_groupi_n_1339 = ((csa_tree_add_69_2_groupi_n_1240 & csa_tree_add_69_2_groupi_n_1176)
    | ((csa_tree_add_69_2_groupi_n_1176 & csa_tree_add_69_2_groupi_n_903) | (csa_tree_add_69_2_groupi_n_903
    & csa_tree_add_69_2_groupi_n_1240)));
 assign csa_tree_add_69_2_groupi_n_1340 = (csa_tree_add_69_2_groupi_n_1176 ^ (csa_tree_add_69_2_groupi_n_903
    ^ csa_tree_add_69_2_groupi_n_1240));
 assign csa_tree_add_69_2_groupi_n_1337 = ((csa_tree_add_69_2_groupi_n_1236 & csa_tree_add_69_2_groupi_n_1118)
    | ((csa_tree_add_69_2_groupi_n_1118 & csa_tree_add_69_2_groupi_n_920) | (csa_tree_add_69_2_groupi_n_920
    & csa_tree_add_69_2_groupi_n_1236)));
 assign csa_tree_add_69_2_groupi_n_1338 = (csa_tree_add_69_2_groupi_n_1118 ^ (csa_tree_add_69_2_groupi_n_920
    ^ csa_tree_add_69_2_groupi_n_1236));
 assign csa_tree_add_69_2_groupi_n_1335 = ((csa_tree_add_69_2_groupi_n_1241 & csa_tree_add_69_2_groupi_n_1114)
    | ((csa_tree_add_69_2_groupi_n_1114 & csa_tree_add_69_2_groupi_n_1177) | (csa_tree_add_69_2_groupi_n_1177
    & csa_tree_add_69_2_groupi_n_1241)));
 assign csa_tree_add_69_2_groupi_n_1336 = (csa_tree_add_69_2_groupi_n_1114 ^ (csa_tree_add_69_2_groupi_n_1177
    ^ csa_tree_add_69_2_groupi_n_1241));
 assign csa_tree_add_69_2_groupi_n_1333 = ((csa_tree_add_69_2_groupi_n_1229 & csa_tree_add_69_2_groupi_n_1100)
    | ((csa_tree_add_69_2_groupi_n_1100 & csa_tree_add_69_2_groupi_n_921) | (csa_tree_add_69_2_groupi_n_921
    & csa_tree_add_69_2_groupi_n_1229)));
 assign csa_tree_add_69_2_groupi_n_1334 = (csa_tree_add_69_2_groupi_n_1100 ^ (csa_tree_add_69_2_groupi_n_921
    ^ csa_tree_add_69_2_groupi_n_1229));
 assign csa_tree_add_69_2_groupi_n_1331 = ((csa_tree_add_69_2_groupi_n_1247 & csa_tree_add_69_2_groupi_n_1124)
    | ((csa_tree_add_69_2_groupi_n_1124 & csa_tree_add_69_2_groupi_n_1158) | (csa_tree_add_69_2_groupi_n_1158
    & csa_tree_add_69_2_groupi_n_1247)));
 assign csa_tree_add_69_2_groupi_n_1332 = (csa_tree_add_69_2_groupi_n_1124 ^ (csa_tree_add_69_2_groupi_n_1158
    ^ csa_tree_add_69_2_groupi_n_1247));
 assign csa_tree_add_69_2_groupi_n_1329 = ((csa_tree_add_69_2_groupi_n_1238 & csa_tree_add_69_2_groupi_n_1102)
    | ((csa_tree_add_69_2_groupi_n_1102 & csa_tree_add_69_2_groupi_n_907) | (csa_tree_add_69_2_groupi_n_907
    & csa_tree_add_69_2_groupi_n_1238)));
 assign csa_tree_add_69_2_groupi_n_1330 = (csa_tree_add_69_2_groupi_n_1102 ^ (csa_tree_add_69_2_groupi_n_907
    ^ csa_tree_add_69_2_groupi_n_1238));
 assign csa_tree_add_69_2_groupi_n_1327 = ((csa_tree_add_69_2_groupi_n_1231 & csa_tree_add_69_2_groupi_n_1106)
    | ((csa_tree_add_69_2_groupi_n_1106 & csa_tree_add_69_2_groupi_n_919) | (csa_tree_add_69_2_groupi_n_919
    & csa_tree_add_69_2_groupi_n_1231)));
 assign csa_tree_add_69_2_groupi_n_1328 = (csa_tree_add_69_2_groupi_n_1106 ^ (csa_tree_add_69_2_groupi_n_919
    ^ csa_tree_add_69_2_groupi_n_1231));
 assign csa_tree_add_69_2_groupi_n_1326 = ((csa_tree_add_69_2_groupi_n_1233 & csa_tree_add_69_2_groupi_n_1088)
    | ((csa_tree_add_69_2_groupi_n_1088 & csa_tree_add_69_2_groupi_n_1085) | (csa_tree_add_69_2_groupi_n_1085
    & csa_tree_add_69_2_groupi_n_1233)));
 assign csa_tree_add_69_2_groupi_n_1357 = (csa_tree_add_69_2_groupi_n_1088 ^ (csa_tree_add_69_2_groupi_n_1085
    ^ csa_tree_add_69_2_groupi_n_1233));
 assign csa_tree_add_69_2_groupi_n_1324 = ((csa_tree_add_69_2_groupi_n_1235 & csa_tree_add_69_2_groupi_n_1134)
    | ((csa_tree_add_69_2_groupi_n_1134 & csa_tree_add_69_2_groupi_n_1185) | (csa_tree_add_69_2_groupi_n_1185
    & csa_tree_add_69_2_groupi_n_1235)));
 assign csa_tree_add_69_2_groupi_n_1325 = (csa_tree_add_69_2_groupi_n_1134 ^ (csa_tree_add_69_2_groupi_n_1185
    ^ csa_tree_add_69_2_groupi_n_1235));
 assign csa_tree_add_69_2_groupi_n_1322 = ((csa_tree_add_69_2_groupi_n_1230 & csa_tree_add_69_2_groupi_n_1164)
    | ((csa_tree_add_69_2_groupi_n_1164 & csa_tree_add_69_2_groupi_n_1101) | (csa_tree_add_69_2_groupi_n_1101
    & csa_tree_add_69_2_groupi_n_1230)));
 assign csa_tree_add_69_2_groupi_n_1323 = (csa_tree_add_69_2_groupi_n_1164 ^ (csa_tree_add_69_2_groupi_n_1101
    ^ csa_tree_add_69_2_groupi_n_1230));
 assign csa_tree_add_69_2_groupi_n_1320 = ((csa_tree_add_69_2_groupi_n_1237 & csa_tree_add_69_2_groupi_n_1116)
    | ((csa_tree_add_69_2_groupi_n_1116 & csa_tree_add_69_2_groupi_n_1119) | (csa_tree_add_69_2_groupi_n_1119
    & csa_tree_add_69_2_groupi_n_1237)));
 assign csa_tree_add_69_2_groupi_n_1321 = (csa_tree_add_69_2_groupi_n_1116 ^ (csa_tree_add_69_2_groupi_n_1119
    ^ csa_tree_add_69_2_groupi_n_1237));
 assign csa_tree_add_69_2_groupi_n_1318 = ((csa_tree_add_69_2_groupi_n_1232 & csa_tree_add_69_2_groupi_n_1120)
    | ((csa_tree_add_69_2_groupi_n_1120 & csa_tree_add_69_2_groupi_n_1107) | (csa_tree_add_69_2_groupi_n_1107
    & csa_tree_add_69_2_groupi_n_1232)));
 assign csa_tree_add_69_2_groupi_n_1319 = (csa_tree_add_69_2_groupi_n_1120 ^ (csa_tree_add_69_2_groupi_n_1107
    ^ csa_tree_add_69_2_groupi_n_1232));
 assign csa_tree_add_69_2_groupi_n_1317 = ~(csa_tree_add_69_2_groupi_n_1312 | csa_tree_add_69_2_groupi_n_1286);
 assign csa_tree_add_69_2_groupi_n_1316 = ~(csa_tree_add_69_2_groupi_n_1312 & csa_tree_add_69_2_groupi_n_1286);
 assign csa_tree_add_69_2_groupi_n_1314 = ~(csa_tree_add_69_2_groupi_n_1289 ^ csa_tree_add_69_2_groupi_n_1297);
 assign csa_tree_add_69_2_groupi_n_1315 = ~(csa_tree_add_69_2_groupi_n_1257 | (csa_tree_add_69_2_groupi_n_1258
    & csa_tree_add_69_2_groupi_n_1254));
 assign csa_tree_add_69_2_groupi_n_1313 = ~(csa_tree_add_69_2_groupi_n_1285 ^ csa_tree_add_69_2_groupi_n_1254);
 assign csa_tree_add_69_2_groupi_n_1312 = ~csa_tree_add_69_2_groupi_n_1301;
 assign csa_tree_add_69_2_groupi_n_1306 = ((csa_tree_add_69_2_groupi_n_1104 & csa_tree_add_69_2_groupi_n_1133)
    | ((csa_tree_add_69_2_groupi_n_1133 & csa_tree_add_69_2_groupi_n_1087) | (csa_tree_add_69_2_groupi_n_1087
    & csa_tree_add_69_2_groupi_n_1104)));
 assign csa_tree_add_69_2_groupi_n_1307 = (csa_tree_add_69_2_groupi_n_1133 ^ (csa_tree_add_69_2_groupi_n_1087
    ^ csa_tree_add_69_2_groupi_n_1104));
 assign csa_tree_add_69_2_groupi_n_1304 = ((csa_tree_add_69_2_groupi_n_1269 & csa_tree_add_69_2_groupi_n_1035)
    | ((csa_tree_add_69_2_groupi_n_1035 & csa_tree_add_69_2_groupi_n_1169) | (csa_tree_add_69_2_groupi_n_1169
    & csa_tree_add_69_2_groupi_n_1269)));
 assign csa_tree_add_69_2_groupi_n_1305 = (csa_tree_add_69_2_groupi_n_1035 ^ (csa_tree_add_69_2_groupi_n_1169
    ^ csa_tree_add_69_2_groupi_n_1269));
 assign csa_tree_add_69_2_groupi_n_1310 = ((csa_tree_add_69_2_groupi_n_1163 & csa_tree_add_69_2_groupi_n_794)
    | ((csa_tree_add_69_2_groupi_n_794 & csa_tree_add_69_2_groupi_n_1095) | (csa_tree_add_69_2_groupi_n_1095
    & csa_tree_add_69_2_groupi_n_1163)));
 assign csa_tree_add_69_2_groupi_n_1311 = (csa_tree_add_69_2_groupi_n_794 ^ (csa_tree_add_69_2_groupi_n_1095
    ^ csa_tree_add_69_2_groupi_n_1163));
 assign csa_tree_add_69_2_groupi_n_1309 = ~(csa_tree_add_69_2_groupi_n_1224 & (csa_tree_add_69_2_groupi_n_1219
    | csa_tree_add_69_2_groupi_n_1223));
 assign csa_tree_add_69_2_groupi_n_1308 = ~((csa_tree_add_69_2_groupi_n_1138 & ~csa_tree_add_69_2_groupi_n_48)
    | (csa_tree_add_69_2_groupi_n_1196 & csa_tree_add_69_2_groupi_n_48));
 assign csa_tree_add_69_2_groupi_n_1303 = ~(csa_tree_add_69_2_groupi_n_1291 ^ csa_tree_add_69_2_groupi_n_1025);
 assign csa_tree_add_69_2_groupi_n_1299 = ((csa_tree_add_69_2_groupi_n_1243 & csa_tree_add_69_2_groupi_n_1043)
    | ((csa_tree_add_69_2_groupi_n_1043 & csa_tree_add_69_2_groupi_n_985) | (csa_tree_add_69_2_groupi_n_985
    & csa_tree_add_69_2_groupi_n_1243)));
 assign csa_tree_add_69_2_groupi_n_1300 = (csa_tree_add_69_2_groupi_n_1043 ^ (csa_tree_add_69_2_groupi_n_985
    ^ csa_tree_add_69_2_groupi_n_1243));
 assign csa_tree_add_69_2_groupi_n_1297 = ((csa_tree_add_69_2_groupi_n_1161 & csa_tree_add_69_2_groupi_n_1147)
    | ((csa_tree_add_69_2_groupi_n_1147 & csa_tree_add_69_2_groupi_n_1137) | (csa_tree_add_69_2_groupi_n_1137
    & csa_tree_add_69_2_groupi_n_1161)));
 assign csa_tree_add_69_2_groupi_n_1298 = (csa_tree_add_69_2_groupi_n_1147 ^ (csa_tree_add_69_2_groupi_n_1137
    ^ csa_tree_add_69_2_groupi_n_1161));
 assign csa_tree_add_69_2_groupi_n_1301 = ~(csa_tree_add_69_2_groupi_n_46 | csa_tree_add_69_2_groupi_n_1206);
 assign csa_tree_add_69_2_groupi_n_1294 = ~(csa_tree_add_69_2_groupi_n_1292 | csa_tree_add_69_2_groupi_n_43);
 assign csa_tree_add_69_2_groupi_n_1293 = ~(csa_tree_add_69_2_groupi_n_1216 ^ csa_tree_add_69_2_groupi_n_1212);
 assign csa_tree_add_69_2_groupi_n_1292 = ~(csa_tree_add_69_2_groupi_n_1094 | ~(csa_tree_add_69_2_groupi_n_1198
    | csa_tree_add_69_2_groupi_n_1011));
 assign csa_tree_add_69_2_groupi_n_1291 = ~((csa_tree_add_69_2_groupi_n_1248 & ~csa_tree_add_69_2_groupi_n_1086)
    | (csa_tree_add_69_2_groupi_n_1249 & csa_tree_add_69_2_groupi_n_1086));
 assign csa_tree_add_69_2_groupi_n_1290 = ~(csa_tree_add_69_2_groupi_n_1222 ^ csa_tree_add_69_2_groupi_n_1076);
 assign csa_tree_add_69_2_groupi_n_1289 = ~(csa_tree_add_69_2_groupi_n_1221 ^ csa_tree_add_69_2_groupi_n_1136);
 assign csa_tree_add_69_2_groupi_n_1285 = ~((csa_tree_add_69_2_groupi_n_1252 & ~csa_tree_add_69_2_groupi_n_1139)
    | (csa_tree_add_69_2_groupi_n_1251 & csa_tree_add_69_2_groupi_n_1139));
 assign csa_tree_add_69_2_groupi_n_1288 = ~(csa_tree_add_69_2_groupi_n_1256 | csa_tree_add_69_2_groupi_n_27);
 assign csa_tree_add_69_2_groupi_n_1284 = ~((csa_tree_add_69_2_groupi_n_1200 & ~csa_tree_add_69_2_groupi_n_1220)
    | (csa_tree_add_69_2_groupi_n_1090 & csa_tree_add_69_2_groupi_n_1220));
 assign csa_tree_add_69_2_groupi_n_1287 = ~(csa_tree_add_69_2_groupi_n_1253 & csa_tree_add_69_2_groupi_n_42);
 assign csa_tree_add_69_2_groupi_n_1286 = ~(csa_tree_add_69_2_groupi_n_1203 ^ csa_tree_add_69_2_groupi_n_1211);
 assign csa_tree_add_69_2_groupi_n_1283 = ~(csa_tree_add_69_2_groupi_n_1208 & (csa_tree_add_69_2_groupi_n_1209
    | csa_tree_add_69_2_groupi_n_1250));
 assign csa_tree_add_69_2_groupi_n_1282 = ~csa_tree_add_69_2_groupi_n_1281;
 assign csa_tree_add_69_2_groupi_n_1280 = ~csa_tree_add_69_2_groupi_n_1218;
 assign csa_tree_add_69_2_groupi_n_1278 = ((csa_tree_add_69_2_groupi_n_1040 & csa_tree_add_69_2_groupi_n_786)
    | ((csa_tree_add_69_2_groupi_n_786 & csa_tree_add_69_2_groupi_n_1037) | (csa_tree_add_69_2_groupi_n_1037
    & csa_tree_add_69_2_groupi_n_1040)));
 assign csa_tree_add_69_2_groupi_n_1279 = (csa_tree_add_69_2_groupi_n_786 ^ (csa_tree_add_69_2_groupi_n_1037
    ^ csa_tree_add_69_2_groupi_n_1040));
 assign csa_tree_add_69_2_groupi_n_1276 = ((csa_tree_add_69_2_groupi_n_1054 & csa_tree_add_69_2_groupi_n_787)
    | ((csa_tree_add_69_2_groupi_n_787 & csa_tree_add_69_2_groupi_n_1063) | (csa_tree_add_69_2_groupi_n_1063
    & csa_tree_add_69_2_groupi_n_1054)));
 assign csa_tree_add_69_2_groupi_n_1277 = (csa_tree_add_69_2_groupi_n_787 ^ (csa_tree_add_69_2_groupi_n_1063
    ^ csa_tree_add_69_2_groupi_n_1054));
 assign csa_tree_add_69_2_groupi_n_1274 = ((csa_tree_add_69_2_groupi_n_1048 & csa_tree_add_69_2_groupi_n_781)
    | ((csa_tree_add_69_2_groupi_n_781 & csa_tree_add_69_2_groupi_n_1039) | (csa_tree_add_69_2_groupi_n_1039
    & csa_tree_add_69_2_groupi_n_1048)));
 assign csa_tree_add_69_2_groupi_n_1275 = (csa_tree_add_69_2_groupi_n_781 ^ (csa_tree_add_69_2_groupi_n_1039
    ^ csa_tree_add_69_2_groupi_n_1048));
 assign csa_tree_add_69_2_groupi_n_1272 = ((csa_tree_add_69_2_groupi_n_1064 & csa_tree_add_69_2_groupi_n_780)
    | ((csa_tree_add_69_2_groupi_n_780 & csa_tree_add_69_2_groupi_n_1041) | (csa_tree_add_69_2_groupi_n_1041
    & csa_tree_add_69_2_groupi_n_1064)));
 assign csa_tree_add_69_2_groupi_n_1273 = (csa_tree_add_69_2_groupi_n_780 ^ (csa_tree_add_69_2_groupi_n_1041
    ^ csa_tree_add_69_2_groupi_n_1064));
 assign csa_tree_add_69_2_groupi_n_1270 = ((csa_tree_add_69_2_groupi_n_1168 & csa_tree_add_69_2_groupi_n_675)
    | ((csa_tree_add_69_2_groupi_n_675 & csa_tree_add_69_2_groupi_n_1044) | (csa_tree_add_69_2_groupi_n_1044
    & csa_tree_add_69_2_groupi_n_1168)));
 assign csa_tree_add_69_2_groupi_n_1271 = (csa_tree_add_69_2_groupi_n_675 ^ (csa_tree_add_69_2_groupi_n_1044
    ^ csa_tree_add_69_2_groupi_n_1168));
 assign csa_tree_add_69_2_groupi_n_1269 = ((csa_tree_add_69_2_groupi_n_39 & csa_tree_add_69_2_groupi_n_890)
    | ((csa_tree_add_69_2_groupi_n_890 & csa_tree_add_69_2_groupi_n_889) | (csa_tree_add_69_2_groupi_n_889
    & csa_tree_add_69_2_groupi_n_39)));
 assign csa_tree_add_69_2_groupi_n_1281 = (csa_tree_add_69_2_groupi_n_890 ^ (csa_tree_add_69_2_groupi_n_889
    ^ csa_tree_add_69_2_groupi_n_39));
 assign csa_tree_add_69_2_groupi_n_1267 = ((csa_tree_add_69_2_groupi_n_1042 & csa_tree_add_69_2_groupi_n_776)
    | ((csa_tree_add_69_2_groupi_n_776 & csa_tree_add_69_2_groupi_n_1067) | (csa_tree_add_69_2_groupi_n_1067
    & csa_tree_add_69_2_groupi_n_1042)));
 assign csa_tree_add_69_2_groupi_n_1268 = (csa_tree_add_69_2_groupi_n_776 ^ (csa_tree_add_69_2_groupi_n_1067
    ^ csa_tree_add_69_2_groupi_n_1042));
 assign csa_tree_add_69_2_groupi_n_1265 = ((csa_tree_add_69_2_groupi_n_1056 & csa_tree_add_69_2_groupi_n_789)
    | ((csa_tree_add_69_2_groupi_n_789 & csa_tree_add_69_2_groupi_n_1029) | (csa_tree_add_69_2_groupi_n_1029
    & csa_tree_add_69_2_groupi_n_1056)));
 assign csa_tree_add_69_2_groupi_n_1266 = (csa_tree_add_69_2_groupi_n_789 ^ (csa_tree_add_69_2_groupi_n_1029
    ^ csa_tree_add_69_2_groupi_n_1056));
 assign csa_tree_add_69_2_groupi_n_1263 = ((csa_tree_add_69_2_groupi_n_1052 & csa_tree_add_69_2_groupi_n_1033)
    | ((csa_tree_add_69_2_groupi_n_1033 & csa_tree_add_69_2_groupi_n_790) | (csa_tree_add_69_2_groupi_n_790
    & csa_tree_add_69_2_groupi_n_1052)));
 assign csa_tree_add_69_2_groupi_n_1264 = (csa_tree_add_69_2_groupi_n_1033 ^ (csa_tree_add_69_2_groupi_n_790
    ^ csa_tree_add_69_2_groupi_n_1052));
 assign csa_tree_add_69_2_groupi_n_1261 = ((csa_tree_add_69_2_groupi_n_1058 & csa_tree_add_69_2_groupi_n_906)
    | ((csa_tree_add_69_2_groupi_n_906 & csa_tree_add_69_2_groupi_n_1065) | (csa_tree_add_69_2_groupi_n_1065
    & csa_tree_add_69_2_groupi_n_1058)));
 assign csa_tree_add_69_2_groupi_n_1262 = (csa_tree_add_69_2_groupi_n_906 ^ (csa_tree_add_69_2_groupi_n_1065
    ^ csa_tree_add_69_2_groupi_n_1058));
 assign csa_tree_add_69_2_groupi_n_1259 = ((csa_tree_add_69_2_groupi_n_1046 & csa_tree_add_69_2_groupi_n_791)
    | ((csa_tree_add_69_2_groupi_n_791 & csa_tree_add_69_2_groupi_n_1061) | (csa_tree_add_69_2_groupi_n_1061
    & csa_tree_add_69_2_groupi_n_1046)));
 assign csa_tree_add_69_2_groupi_n_1260 = (csa_tree_add_69_2_groupi_n_791 ^ (csa_tree_add_69_2_groupi_n_1061
    ^ csa_tree_add_69_2_groupi_n_1046));
 assign csa_tree_add_69_2_groupi_n_1258 = ~(csa_tree_add_69_2_groupi_n_1197 & ~csa_tree_add_69_2_groupi_n_1252);
 assign csa_tree_add_69_2_groupi_n_1257 = ~(csa_tree_add_69_2_groupi_n_1197 | ~csa_tree_add_69_2_groupi_n_1252);
 assign csa_tree_add_69_2_groupi_n_1256 = ~(csa_tree_add_69_2_groupi_n_1144 | ~csa_tree_add_69_2_groupi_n_1211);
 assign csa_tree_add_69_2_groupi_n_1253 = ~(csa_tree_add_69_2_groupi_n_40 & ~csa_tree_add_69_2_groupi_n_1249);
 assign csa_tree_add_69_2_groupi_n_1255 = ~(csa_tree_add_69_2_groupi_n_1194 ^ csa_tree_add_69_2_groupi_n_1213);
 assign csa_tree_add_69_2_groupi_n_1254 = ~(csa_tree_add_69_2_groupi_n_1210 & (csa_tree_add_69_2_groupi_n_1207
    | csa_tree_add_69_2_groupi_n_1141));
 assign csa_tree_add_69_2_groupi_n_1252 = ~csa_tree_add_69_2_groupi_n_1251;
 assign csa_tree_add_69_2_groupi_n_1249 = ~csa_tree_add_69_2_groupi_n_1248;
 assign csa_tree_add_69_2_groupi_n_1246 = ((csa_tree_add_69_2_groupi_n_1027 & csa_tree_add_69_2_groupi_n_796)
    | ((csa_tree_add_69_2_groupi_n_796 & csa_tree_add_69_2_groupi_n_1068) | (csa_tree_add_69_2_groupi_n_1068
    & csa_tree_add_69_2_groupi_n_1027)));
 assign csa_tree_add_69_2_groupi_n_1247 = (csa_tree_add_69_2_groupi_n_796 ^ (csa_tree_add_69_2_groupi_n_1068
    ^ csa_tree_add_69_2_groupi_n_1027));
 assign csa_tree_add_69_2_groupi_n_1244 = ((csa_tree_add_69_2_groupi_n_1059 & csa_tree_add_69_2_groupi_n_778)
    | ((csa_tree_add_69_2_groupi_n_778 & csa_tree_add_69_2_groupi_n_1070) | (csa_tree_add_69_2_groupi_n_1070
    & csa_tree_add_69_2_groupi_n_1059)));
 assign csa_tree_add_69_2_groupi_n_1245 = (csa_tree_add_69_2_groupi_n_778 ^ (csa_tree_add_69_2_groupi_n_1070
    ^ csa_tree_add_69_2_groupi_n_1059));
 assign csa_tree_add_69_2_groupi_n_1242 = ((csa_tree_add_69_2_groupi_n_1060 & csa_tree_add_69_2_groupi_n_784)
    | ((csa_tree_add_69_2_groupi_n_784 & csa_tree_add_69_2_groupi_n_807) | (csa_tree_add_69_2_groupi_n_807
    & csa_tree_add_69_2_groupi_n_1060)));
 assign csa_tree_add_69_2_groupi_n_1243 = (csa_tree_add_69_2_groupi_n_784 ^ (csa_tree_add_69_2_groupi_n_807
    ^ csa_tree_add_69_2_groupi_n_1060));
 assign csa_tree_add_69_2_groupi_n_1240 = ((csa_tree_add_69_2_groupi_n_1031 & csa_tree_add_69_2_groupi_n_774)
    | ((csa_tree_add_69_2_groupi_n_774 & csa_tree_add_69_2_groupi_n_1062) | (csa_tree_add_69_2_groupi_n_1062
    & csa_tree_add_69_2_groupi_n_1031)));
 assign csa_tree_add_69_2_groupi_n_1241 = (csa_tree_add_69_2_groupi_n_774 ^ (csa_tree_add_69_2_groupi_n_1062
    ^ csa_tree_add_69_2_groupi_n_1031));
 assign csa_tree_add_69_2_groupi_n_1250 = ((csa_tree_add_69_2_groupi_n_995 & csa_tree_add_69_2_groupi_n_835)
    | ((csa_tree_add_69_2_groupi_n_835 & csa_tree_add_69_2_groupi_n_834) | (csa_tree_add_69_2_groupi_n_834
    & csa_tree_add_69_2_groupi_n_995)));
 assign csa_tree_add_69_2_groupi_n_1251 = (csa_tree_add_69_2_groupi_n_835 ^ (csa_tree_add_69_2_groupi_n_834
    ^ csa_tree_add_69_2_groupi_n_995));
 assign csa_tree_add_69_2_groupi_n_1238 = ((csa_tree_add_69_2_groupi_n_1045 & csa_tree_add_69_2_groupi_n_785)
    | ((csa_tree_add_69_2_groupi_n_785 & csa_tree_add_69_2_groupi_n_1038) | (csa_tree_add_69_2_groupi_n_1038
    & csa_tree_add_69_2_groupi_n_1045)));
 assign csa_tree_add_69_2_groupi_n_1239 = (csa_tree_add_69_2_groupi_n_785 ^ (csa_tree_add_69_2_groupi_n_1038
    ^ csa_tree_add_69_2_groupi_n_1045));
 assign csa_tree_add_69_2_groupi_n_1236 = ((csa_tree_add_69_2_groupi_n_1055 & csa_tree_add_69_2_groupi_n_793)
    | ((csa_tree_add_69_2_groupi_n_793 & csa_tree_add_69_2_groupi_n_1032) | (csa_tree_add_69_2_groupi_n_1032
    & csa_tree_add_69_2_groupi_n_1055)));
 assign csa_tree_add_69_2_groupi_n_1237 = (csa_tree_add_69_2_groupi_n_793 ^ (csa_tree_add_69_2_groupi_n_1032
    ^ csa_tree_add_69_2_groupi_n_1055));
 assign csa_tree_add_69_2_groupi_n_1234 = ((csa_tree_add_69_2_groupi_n_1047 & csa_tree_add_69_2_groupi_n_925)
    | ((csa_tree_add_69_2_groupi_n_925 & csa_tree_add_69_2_groupi_n_1066) | (csa_tree_add_69_2_groupi_n_1066
    & csa_tree_add_69_2_groupi_n_1047)));
 assign csa_tree_add_69_2_groupi_n_1235 = (csa_tree_add_69_2_groupi_n_925 ^ (csa_tree_add_69_2_groupi_n_1066
    ^ csa_tree_add_69_2_groupi_n_1047));
 assign csa_tree_add_69_2_groupi_n_1233 = ((csa_tree_add_69_2_groupi_n_1036 & csa_tree_add_69_2_groupi_n_830)
    | ((csa_tree_add_69_2_groupi_n_830 & csa_tree_add_69_2_groupi_n_811) | (csa_tree_add_69_2_groupi_n_811
    & csa_tree_add_69_2_groupi_n_1036)));
 assign csa_tree_add_69_2_groupi_n_1248 = (csa_tree_add_69_2_groupi_n_830 ^ (csa_tree_add_69_2_groupi_n_811
    ^ csa_tree_add_69_2_groupi_n_1036));
 assign csa_tree_add_69_2_groupi_n_1231 = ((csa_tree_add_69_2_groupi_n_1051 & csa_tree_add_69_2_groupi_n_792)
    | ((csa_tree_add_69_2_groupi_n_792 & csa_tree_add_69_2_groupi_n_1050) | (csa_tree_add_69_2_groupi_n_1050
    & csa_tree_add_69_2_groupi_n_1051)));
 assign csa_tree_add_69_2_groupi_n_1232 = (csa_tree_add_69_2_groupi_n_792 ^ (csa_tree_add_69_2_groupi_n_1050
    ^ csa_tree_add_69_2_groupi_n_1051));
 assign csa_tree_add_69_2_groupi_n_1229 = ((csa_tree_add_69_2_groupi_n_1049 & csa_tree_add_69_2_groupi_n_795)
    | ((csa_tree_add_69_2_groupi_n_795 & csa_tree_add_69_2_groupi_n_1028) | (csa_tree_add_69_2_groupi_n_1028
    & csa_tree_add_69_2_groupi_n_1049)));
 assign csa_tree_add_69_2_groupi_n_1230 = (csa_tree_add_69_2_groupi_n_795 ^ (csa_tree_add_69_2_groupi_n_1028
    ^ csa_tree_add_69_2_groupi_n_1049));
 assign csa_tree_add_69_2_groupi_n_1227 = ((csa_tree_add_69_2_groupi_n_1053 & csa_tree_add_69_2_groupi_n_783)
    | ((csa_tree_add_69_2_groupi_n_783 & csa_tree_add_69_2_groupi_n_1030) | (csa_tree_add_69_2_groupi_n_1030
    & csa_tree_add_69_2_groupi_n_1053)));
 assign csa_tree_add_69_2_groupi_n_1228 = (csa_tree_add_69_2_groupi_n_783 ^ (csa_tree_add_69_2_groupi_n_1030
    ^ csa_tree_add_69_2_groupi_n_1053));
 assign csa_tree_add_69_2_groupi_n_1225 = ((csa_tree_add_69_2_groupi_n_1069 & csa_tree_add_69_2_groupi_n_788)
    | ((csa_tree_add_69_2_groupi_n_788 & csa_tree_add_69_2_groupi_n_1034) | (csa_tree_add_69_2_groupi_n_1034
    & csa_tree_add_69_2_groupi_n_1069)));
 assign csa_tree_add_69_2_groupi_n_1226 = (csa_tree_add_69_2_groupi_n_788 ^ (csa_tree_add_69_2_groupi_n_1034
    ^ csa_tree_add_69_2_groupi_n_1069));
 assign csa_tree_add_69_2_groupi_n_1224 = ~(csa_tree_add_69_2_groupi_n_1195 & csa_tree_add_69_2_groupi_n_1213);
 assign csa_tree_add_69_2_groupi_n_1223 = ~(csa_tree_add_69_2_groupi_n_1195 | csa_tree_add_69_2_groupi_n_1213);
 assign csa_tree_add_69_2_groupi_n_1222 = ~(csa_tree_add_69_2_groupi_n_731 ^ csa_tree_add_69_2_groupi_n_1153);
 assign csa_tree_add_69_2_groupi_n_1221 = ~(csa_tree_add_69_2_groupi_n_1149 ^ csa_tree_add_69_2_groupi_n_1097);
 assign csa_tree_add_69_2_groupi_n_1220 = ~((csa_tree_add_69_2_groupi_n_1140 & ~csa_tree_add_69_2_groupi_n_1141)
    | (csa_tree_add_69_2_groupi_n_1199 & csa_tree_add_69_2_groupi_n_1141));
 assign csa_tree_add_69_2_groupi_n_1217 = ~(csa_tree_add_69_2_groupi_n_1198 ^ csa_tree_add_69_2_groupi_n_1011);
 assign csa_tree_add_69_2_groupi_n_1216 = ~((csa_tree_add_69_2_groupi_n_1193 & ~n_447) | (csa_tree_add_69_2_groupi_n_1192
    & n_447));
 assign csa_tree_add_69_2_groupi_n_1219 = ~(csa_tree_add_69_2_groupi_n_994 ^ (csa_tree_add_69_2_groupi_n_862
    ^ csa_tree_add_69_2_groupi_n_1142));
 assign csa_tree_add_69_2_groupi_n_1218 = ~(csa_tree_add_69_2_groupi_n_1205 | csa_tree_add_69_2_groupi_n_37);
 assign csa_tree_add_69_2_groupi_n_1215 = ~(csa_tree_add_69_2_groupi_n_45 & csa_tree_add_69_2_groupi_n_36);
 assign csa_tree_add_69_2_groupi_n_1213 = ((csa_tree_add_69_2_groupi_n_854 & csa_tree_add_69_2_groupi_n_1003)
    | ((csa_tree_add_69_2_groupi_n_1003 & csa_tree_add_69_2_groupi_n_663) | (csa_tree_add_69_2_groupi_n_663
    & csa_tree_add_69_2_groupi_n_854)));
 assign csa_tree_add_69_2_groupi_n_1214 = (csa_tree_add_69_2_groupi_n_1003 ^ (csa_tree_add_69_2_groupi_n_663
    ^ csa_tree_add_69_2_groupi_n_854));
 assign csa_tree_add_69_2_groupi_n_1211 = ((csa_tree_add_69_2_groupi_n_942 & csa_tree_add_69_2_groupi_n_893)
    | ((csa_tree_add_69_2_groupi_n_893 & csa_tree_add_69_2_groupi_n_777) | (csa_tree_add_69_2_groupi_n_777
    & csa_tree_add_69_2_groupi_n_942)));
 assign csa_tree_add_69_2_groupi_n_1212 = (csa_tree_add_69_2_groupi_n_893 ^ (csa_tree_add_69_2_groupi_n_777
    ^ csa_tree_add_69_2_groupi_n_942));
 assign csa_tree_add_69_2_groupi_n_1210 = ~(csa_tree_add_69_2_groupi_n_1200 & ~csa_tree_add_69_2_groupi_n_1140);
 assign csa_tree_add_69_2_groupi_n_1209 = ~(csa_tree_add_69_2_groupi_n_1202 | csa_tree_add_69_2_groupi_n_1196);
 assign csa_tree_add_69_2_groupi_n_1208 = ~(csa_tree_add_69_2_groupi_n_1202 & csa_tree_add_69_2_groupi_n_1196);
 assign csa_tree_add_69_2_groupi_n_1207 = ~(csa_tree_add_69_2_groupi_n_1200 | csa_tree_add_69_2_groupi_n_1199);
 assign csa_tree_add_69_2_groupi_n_1206 = ~(n_447 | csa_tree_add_69_2_groupi_n_1193);
 assign csa_tree_add_69_2_groupi_n_1205 = ~(csa_tree_add_69_2_groupi_n_1084 | csa_tree_add_69_2_groupi_n_1093);
 assign csa_tree_add_69_2_groupi_n_1203 = ~((csa_tree_add_69_2_groupi_n_1024 & ~csa_tree_add_69_2_groupi_n_865)
    | (csa_tree_add_69_2_groupi_n_1143 & csa_tree_add_69_2_groupi_n_865));
 assign csa_tree_add_69_2_groupi_n_1202 = ~csa_tree_add_69_2_groupi_n_1091;
 assign csa_tree_add_69_2_groupi_n_1201 = ~csa_tree_add_69_2_groupi_n_1092;
 assign csa_tree_add_69_2_groupi_n_1200 = ~csa_tree_add_69_2_groupi_n_1090;
 assign csa_tree_add_69_2_groupi_n_1199 = ~csa_tree_add_69_2_groupi_n_1140;
 assign csa_tree_add_69_2_groupi_n_1197 = ~csa_tree_add_69_2_groupi_n_1139;
 assign csa_tree_add_69_2_groupi_n_1196 = ~csa_tree_add_69_2_groupi_n_1138;
 assign csa_tree_add_69_2_groupi_n_1195 = ~csa_tree_add_69_2_groupi_n_1194;
 assign csa_tree_add_69_2_groupi_n_1192 = ~csa_tree_add_69_2_groupi_n_1193;
 assign csa_tree_add_69_2_groupi_n_1190 = ((csa_tree_add_69_2_groupi_n_727 & csa_tree_add_69_2_groupi_n_658)
    | ((csa_tree_add_69_2_groupi_n_658 & csa_tree_add_69_2_groupi_n_901) | (csa_tree_add_69_2_groupi_n_901
    & csa_tree_add_69_2_groupi_n_727)));
 assign csa_tree_add_69_2_groupi_n_1191 = (csa_tree_add_69_2_groupi_n_658 ^ (csa_tree_add_69_2_groupi_n_901
    ^ csa_tree_add_69_2_groupi_n_727));
 assign csa_tree_add_69_2_groupi_n_1188 = ((csa_tree_add_69_2_groupi_n_839 & csa_tree_add_69_2_groupi_n_826)
    | ((csa_tree_add_69_2_groupi_n_826 & csa_tree_add_69_2_groupi_n_805) | (csa_tree_add_69_2_groupi_n_805
    & csa_tree_add_69_2_groupi_n_839)));
 assign csa_tree_add_69_2_groupi_n_1189 = (csa_tree_add_69_2_groupi_n_826 ^ (csa_tree_add_69_2_groupi_n_805
    ^ csa_tree_add_69_2_groupi_n_839));
 assign csa_tree_add_69_2_groupi_n_1186 = ((csa_tree_add_69_2_groupi_n_689 & csa_tree_add_69_2_groupi_n_670)
    | ((csa_tree_add_69_2_groupi_n_670 & csa_tree_add_69_2_groupi_n_886) | (csa_tree_add_69_2_groupi_n_886
    & csa_tree_add_69_2_groupi_n_689)));
 assign csa_tree_add_69_2_groupi_n_1187 = (csa_tree_add_69_2_groupi_n_670 ^ (csa_tree_add_69_2_groupi_n_886
    ^ csa_tree_add_69_2_groupi_n_689));
 assign csa_tree_add_69_2_groupi_n_1184 = ((csa_tree_add_69_2_groupi_n_841 & csa_tree_add_69_2_groupi_n_782)
    | ((csa_tree_add_69_2_groupi_n_782 & csa_tree_add_69_2_groupi_n_881) | (csa_tree_add_69_2_groupi_n_881
    & csa_tree_add_69_2_groupi_n_841)));
 assign csa_tree_add_69_2_groupi_n_1185 = (csa_tree_add_69_2_groupi_n_782 ^ (csa_tree_add_69_2_groupi_n_881
    ^ csa_tree_add_69_2_groupi_n_841));
 assign csa_tree_add_69_2_groupi_n_1182 = ((csa_tree_add_69_2_groupi_n_849 & csa_tree_add_69_2_groupi_n_831)
    | ((csa_tree_add_69_2_groupi_n_831 & csa_tree_add_69_2_groupi_n_802) | (csa_tree_add_69_2_groupi_n_802
    & csa_tree_add_69_2_groupi_n_849)));
 assign csa_tree_add_69_2_groupi_n_1183 = (csa_tree_add_69_2_groupi_n_831 ^ (csa_tree_add_69_2_groupi_n_802
    ^ csa_tree_add_69_2_groupi_n_849));
 assign csa_tree_add_69_2_groupi_n_1180 = ((csa_tree_add_69_2_groupi_n_851 & csa_tree_add_69_2_groupi_n_809)
    | ((csa_tree_add_69_2_groupi_n_809 & csa_tree_add_69_2_groupi_n_815) | (csa_tree_add_69_2_groupi_n_815
    & csa_tree_add_69_2_groupi_n_851)));
 assign csa_tree_add_69_2_groupi_n_1181 = (csa_tree_add_69_2_groupi_n_809 ^ (csa_tree_add_69_2_groupi_n_815
    ^ csa_tree_add_69_2_groupi_n_851));
 assign csa_tree_add_69_2_groupi_n_1178 = ((csa_tree_add_69_2_groupi_n_700 & csa_tree_add_69_2_groupi_n_665)
    | ((csa_tree_add_69_2_groupi_n_665 & csa_tree_add_69_2_groupi_n_891) | (csa_tree_add_69_2_groupi_n_891
    & csa_tree_add_69_2_groupi_n_700)));
 assign csa_tree_add_69_2_groupi_n_1179 = (csa_tree_add_69_2_groupi_n_665 ^ (csa_tree_add_69_2_groupi_n_891
    ^ csa_tree_add_69_2_groupi_n_700));
 assign csa_tree_add_69_2_groupi_n_1176 = ((csa_tree_add_69_2_groupi_n_850 & csa_tree_add_69_2_groupi_n_806)
    | ((csa_tree_add_69_2_groupi_n_806 & csa_tree_add_69_2_groupi_n_797) | (csa_tree_add_69_2_groupi_n_797
    & csa_tree_add_69_2_groupi_n_850)));
 assign csa_tree_add_69_2_groupi_n_1177 = (csa_tree_add_69_2_groupi_n_806 ^ (csa_tree_add_69_2_groupi_n_797
    ^ csa_tree_add_69_2_groupi_n_850));
 assign csa_tree_add_69_2_groupi_n_1174 = ((csa_tree_add_69_2_groupi_n_704 & csa_tree_add_69_2_groupi_n_656)
    | ((csa_tree_add_69_2_groupi_n_656 & csa_tree_add_69_2_groupi_n_908) | (csa_tree_add_69_2_groupi_n_908
    & csa_tree_add_69_2_groupi_n_704)));
 assign csa_tree_add_69_2_groupi_n_1175 = (csa_tree_add_69_2_groupi_n_656 ^ (csa_tree_add_69_2_groupi_n_908
    ^ csa_tree_add_69_2_groupi_n_704));
 assign csa_tree_add_69_2_groupi_n_1172 = ((csa_tree_add_69_2_groupi_n_728 & csa_tree_add_69_2_groupi_n_725)
    | ((csa_tree_add_69_2_groupi_n_725 & csa_tree_add_69_2_groupi_n_899) | (csa_tree_add_69_2_groupi_n_899
    & csa_tree_add_69_2_groupi_n_728)));
 assign csa_tree_add_69_2_groupi_n_1173 = (csa_tree_add_69_2_groupi_n_725 ^ (csa_tree_add_69_2_groupi_n_899
    ^ csa_tree_add_69_2_groupi_n_728));
 assign csa_tree_add_69_2_groupi_n_1170 = ((csa_tree_add_69_2_groupi_n_845 & csa_tree_add_69_2_groupi_n_825)
    | ((csa_tree_add_69_2_groupi_n_825 & csa_tree_add_69_2_groupi_n_812) | (csa_tree_add_69_2_groupi_n_812
    & csa_tree_add_69_2_groupi_n_845)));
 assign csa_tree_add_69_2_groupi_n_1171 = (csa_tree_add_69_2_groupi_n_825 ^ (csa_tree_add_69_2_groupi_n_812
    ^ csa_tree_add_69_2_groupi_n_845));
 assign csa_tree_add_69_2_groupi_n_1168 = ((n_450 & csa_tree_add_69_2_groupi_n_775) | ((csa_tree_add_69_2_groupi_n_775
    & csa_tree_add_69_2_groupi_n_804) | (csa_tree_add_69_2_groupi_n_804 & n_450)));
 assign csa_tree_add_69_2_groupi_n_1169 = (csa_tree_add_69_2_groupi_n_775 ^ (csa_tree_add_69_2_groupi_n_804
    ^ n_450));
 assign csa_tree_add_69_2_groupi_n_1166 = ((csa_tree_add_69_2_groupi_n_844 & csa_tree_add_69_2_groupi_n_816)
    | ((csa_tree_add_69_2_groupi_n_816 & csa_tree_add_69_2_groupi_n_813) | (csa_tree_add_69_2_groupi_n_813
    & csa_tree_add_69_2_groupi_n_844)));
 assign csa_tree_add_69_2_groupi_n_1167 = (csa_tree_add_69_2_groupi_n_816 ^ (csa_tree_add_69_2_groupi_n_813
    ^ csa_tree_add_69_2_groupi_n_844));
 assign csa_tree_add_69_2_groupi_n_1164 = ((csa_tree_add_69_2_groupi_n_729 & csa_tree_add_69_2_groupi_n_722)
    | ((csa_tree_add_69_2_groupi_n_722 & csa_tree_add_69_2_groupi_n_916) | (csa_tree_add_69_2_groupi_n_916
    & csa_tree_add_69_2_groupi_n_729)));
 assign csa_tree_add_69_2_groupi_n_1165 = (csa_tree_add_69_2_groupi_n_722 ^ (csa_tree_add_69_2_groupi_n_916
    ^ csa_tree_add_69_2_groupi_n_729));
 assign csa_tree_add_69_2_groupi_n_1163 = ((csa_tree_add_69_2_groupi_n_1004 & csa_tree_add_69_2_groupi_n_662)
    | ((csa_tree_add_69_2_groupi_n_662 & csa_tree_add_69_2_groupi_n_923) | (csa_tree_add_69_2_groupi_n_923
    & csa_tree_add_69_2_groupi_n_1004)));
 assign csa_tree_add_69_2_groupi_n_1198 = (csa_tree_add_69_2_groupi_n_662 ^ (csa_tree_add_69_2_groupi_n_923
    ^ csa_tree_add_69_2_groupi_n_1004));
 assign csa_tree_add_69_2_groupi_n_1193 = ((csa_tree_add_69_2_groupi_n_855 & csa_tree_add_69_2_groupi_n_614)
    | ((csa_tree_add_69_2_groupi_n_614 & csa_tree_add_69_2_groupi_n_924) | (csa_tree_add_69_2_groupi_n_924
    & csa_tree_add_69_2_groupi_n_855)));
 assign csa_tree_add_69_2_groupi_n_1194 = (csa_tree_add_69_2_groupi_n_614 ^ (csa_tree_add_69_2_groupi_n_924
    ^ csa_tree_add_69_2_groupi_n_855));
 assign csa_tree_add_69_2_groupi_n_1161 = ((csa_tree_add_69_2_groupi_n_846 & csa_tree_add_69_2_groupi_n_824)
    | ((csa_tree_add_69_2_groupi_n_824 & csa_tree_add_69_2_groupi_n_911) | (csa_tree_add_69_2_groupi_n_911
    & csa_tree_add_69_2_groupi_n_846)));
 assign csa_tree_add_69_2_groupi_n_1162 = (csa_tree_add_69_2_groupi_n_824 ^ (csa_tree_add_69_2_groupi_n_911
    ^ csa_tree_add_69_2_groupi_n_846));
 assign csa_tree_add_69_2_groupi_n_1159 = ((csa_tree_add_69_2_groupi_n_836 & csa_tree_add_69_2_groupi_n_833)
    | ((csa_tree_add_69_2_groupi_n_833 & csa_tree_add_69_2_groupi_n_801) | (csa_tree_add_69_2_groupi_n_801
    & csa_tree_add_69_2_groupi_n_836)));
 assign csa_tree_add_69_2_groupi_n_1160 = (csa_tree_add_69_2_groupi_n_833 ^ (csa_tree_add_69_2_groupi_n_801
    ^ csa_tree_add_69_2_groupi_n_836));
 assign csa_tree_add_69_2_groupi_n_1157 = ((csa_tree_add_69_2_groupi_n_843 & csa_tree_add_69_2_groupi_n_822)
    | ((csa_tree_add_69_2_groupi_n_822 & csa_tree_add_69_2_groupi_n_819) | (csa_tree_add_69_2_groupi_n_819
    & csa_tree_add_69_2_groupi_n_843)));
 assign csa_tree_add_69_2_groupi_n_1158 = (csa_tree_add_69_2_groupi_n_822 ^ (csa_tree_add_69_2_groupi_n_819
    ^ csa_tree_add_69_2_groupi_n_843));
 assign csa_tree_add_69_2_groupi_n_1155 = ((csa_tree_add_69_2_groupi_n_693 & csa_tree_add_69_2_groupi_n_666)
    | ((csa_tree_add_69_2_groupi_n_666 & csa_tree_add_69_2_groupi_n_896) | (csa_tree_add_69_2_groupi_n_896
    & csa_tree_add_69_2_groupi_n_693)));
 assign csa_tree_add_69_2_groupi_n_1156 = (csa_tree_add_69_2_groupi_n_666 ^ (csa_tree_add_69_2_groupi_n_896
    ^ csa_tree_add_69_2_groupi_n_693));
 assign csa_tree_add_69_2_groupi_n_1153 = ((csa_tree_add_69_2_groupi_n_1057 & csa_tree_add_69_2_groupi_n_909)
    | ((csa_tree_add_69_2_groupi_n_909 & csa_tree_add_69_2_groupi_n_898) | (csa_tree_add_69_2_groupi_n_898
    & csa_tree_add_69_2_groupi_n_1057)));
 assign csa_tree_add_69_2_groupi_n_1154 = (csa_tree_add_69_2_groupi_n_909 ^ (csa_tree_add_69_2_groupi_n_898
    ^ csa_tree_add_69_2_groupi_n_1057));
 assign csa_tree_add_69_2_groupi_n_1151 = ((csa_tree_add_69_2_groupi_n_848 & csa_tree_add_69_2_groupi_n_820)
    | ((csa_tree_add_69_2_groupi_n_820 & csa_tree_add_69_2_groupi_n_800) | (csa_tree_add_69_2_groupi_n_800
    & csa_tree_add_69_2_groupi_n_848)));
 assign csa_tree_add_69_2_groupi_n_1152 = (csa_tree_add_69_2_groupi_n_820 ^ (csa_tree_add_69_2_groupi_n_800
    ^ csa_tree_add_69_2_groupi_n_848));
 assign csa_tree_add_69_2_groupi_n_1149 = ((csa_tree_add_69_2_groupi_n_1015 & csa_tree_add_69_2_groupi_n_721)
    | ((csa_tree_add_69_2_groupi_n_721 & csa_tree_add_69_2_groupi_n_922) | (csa_tree_add_69_2_groupi_n_922
    & csa_tree_add_69_2_groupi_n_1015)));
 assign csa_tree_add_69_2_groupi_n_1150 = (csa_tree_add_69_2_groupi_n_721 ^ (csa_tree_add_69_2_groupi_n_922
    ^ csa_tree_add_69_2_groupi_n_1015));
 assign csa_tree_add_69_2_groupi_n_1147 = ((csa_tree_add_69_2_groupi_n_695 & csa_tree_add_69_2_groupi_n_726)
    | ((csa_tree_add_69_2_groupi_n_726 & csa_tree_add_69_2_groupi_n_904) | (csa_tree_add_69_2_groupi_n_904
    & csa_tree_add_69_2_groupi_n_695)));
 assign csa_tree_add_69_2_groupi_n_1148 = (csa_tree_add_69_2_groupi_n_726 ^ (csa_tree_add_69_2_groupi_n_904
    ^ csa_tree_add_69_2_groupi_n_695));
 assign csa_tree_add_69_2_groupi_n_1145 = ((csa_tree_add_69_2_groupi_n_838 & csa_tree_add_69_2_groupi_n_829)
    | ((csa_tree_add_69_2_groupi_n_829 & csa_tree_add_69_2_groupi_n_808) | (csa_tree_add_69_2_groupi_n_808
    & csa_tree_add_69_2_groupi_n_838)));
 assign csa_tree_add_69_2_groupi_n_1146 = (csa_tree_add_69_2_groupi_n_829 ^ (csa_tree_add_69_2_groupi_n_808
    ^ csa_tree_add_69_2_groupi_n_838));
 assign csa_tree_add_69_2_groupi_n_1144 = ~(csa_tree_add_69_2_groupi_n_1024 | csa_tree_add_69_2_groupi_n_865);
 assign csa_tree_add_69_2_groupi_n_1143 = ~csa_tree_add_69_2_groupi_n_1024;
 assign csa_tree_add_69_2_groupi_n_1136 = ((csa_tree_add_69_2_groupi_n_939 & csa_tree_add_69_2_groupi_n_672)
    | ((csa_tree_add_69_2_groupi_n_672 & csa_tree_add_69_2_groupi_n_884) | (csa_tree_add_69_2_groupi_n_884
    & csa_tree_add_69_2_groupi_n_939)));
 assign csa_tree_add_69_2_groupi_n_1137 = (csa_tree_add_69_2_groupi_n_672 ^ (csa_tree_add_69_2_groupi_n_884
    ^ csa_tree_add_69_2_groupi_n_939));
 assign csa_tree_add_69_2_groupi_n_1134 = ((csa_tree_add_69_2_groupi_n_933 & csa_tree_add_69_2_groupi_n_655)
    | ((csa_tree_add_69_2_groupi_n_655 & csa_tree_add_69_2_groupi_n_717) | (csa_tree_add_69_2_groupi_n_717
    & csa_tree_add_69_2_groupi_n_933)));
 assign csa_tree_add_69_2_groupi_n_1135 = (csa_tree_add_69_2_groupi_n_655 ^ (csa_tree_add_69_2_groupi_n_717
    ^ csa_tree_add_69_2_groupi_n_933));
 assign csa_tree_add_69_2_groupi_n_1132 = ((csa_tree_add_69_2_groupi_n_853 & csa_tree_add_69_2_groupi_n_828)
    | ((csa_tree_add_69_2_groupi_n_828 & csa_tree_add_69_2_groupi_n_823) | (csa_tree_add_69_2_groupi_n_823
    & csa_tree_add_69_2_groupi_n_853)));
 assign csa_tree_add_69_2_groupi_n_1133 = (csa_tree_add_69_2_groupi_n_828 ^ (csa_tree_add_69_2_groupi_n_823
    ^ csa_tree_add_69_2_groupi_n_853));
 assign csa_tree_add_69_2_groupi_n_1130 = ((csa_tree_add_69_2_groupi_n_847 & csa_tree_add_69_2_groupi_n_821)
    | ((csa_tree_add_69_2_groupi_n_821 & csa_tree_add_69_2_groupi_n_814) | (csa_tree_add_69_2_groupi_n_814
    & csa_tree_add_69_2_groupi_n_847)));
 assign csa_tree_add_69_2_groupi_n_1131 = (csa_tree_add_69_2_groupi_n_821 ^ (csa_tree_add_69_2_groupi_n_814
    ^ csa_tree_add_69_2_groupi_n_847));
 assign csa_tree_add_69_2_groupi_n_1128 = ((csa_tree_add_69_2_groupi_n_694 & csa_tree_add_69_2_groupi_n_664)
    | ((csa_tree_add_69_2_groupi_n_664 & csa_tree_add_69_2_groupi_n_897) | (csa_tree_add_69_2_groupi_n_897
    & csa_tree_add_69_2_groupi_n_694)));
 assign csa_tree_add_69_2_groupi_n_1129 = (csa_tree_add_69_2_groupi_n_664 ^ (csa_tree_add_69_2_groupi_n_897
    ^ csa_tree_add_69_2_groupi_n_694));
 assign csa_tree_add_69_2_groupi_n_1126 = ((csa_tree_add_69_2_groupi_n_859 & csa_tree_add_69_2_groupi_n_674)
    | ((csa_tree_add_69_2_groupi_n_674 & csa_tree_add_69_2_groupi_n_668) | (csa_tree_add_69_2_groupi_n_668
    & csa_tree_add_69_2_groupi_n_859)));
 assign csa_tree_add_69_2_groupi_n_1127 = (csa_tree_add_69_2_groupi_n_674 ^ (csa_tree_add_69_2_groupi_n_668
    ^ csa_tree_add_69_2_groupi_n_859));
 assign csa_tree_add_69_2_groupi_n_1124 = ((csa_tree_add_69_2_groupi_n_934 & csa_tree_add_69_2_groupi_n_661)
    | ((csa_tree_add_69_2_groupi_n_661 & csa_tree_add_69_2_groupi_n_723) | (csa_tree_add_69_2_groupi_n_723
    & csa_tree_add_69_2_groupi_n_934)));
 assign csa_tree_add_69_2_groupi_n_1125 = (csa_tree_add_69_2_groupi_n_661 ^ (csa_tree_add_69_2_groupi_n_723
    ^ csa_tree_add_69_2_groupi_n_934));
 assign csa_tree_add_69_2_groupi_n_1122 = ((csa_tree_add_69_2_groupi_n_707 & csa_tree_add_69_2_groupi_n_719)
    | ((csa_tree_add_69_2_groupi_n_719 & csa_tree_add_69_2_groupi_n_913) | (csa_tree_add_69_2_groupi_n_913
    & csa_tree_add_69_2_groupi_n_707)));
 assign csa_tree_add_69_2_groupi_n_1123 = (csa_tree_add_69_2_groupi_n_719 ^ (csa_tree_add_69_2_groupi_n_913
    ^ csa_tree_add_69_2_groupi_n_707));
 assign csa_tree_add_69_2_groupi_n_1120 = ((csa_tree_add_69_2_groupi_n_932 & csa_tree_add_69_2_groupi_n_676)
    | ((csa_tree_add_69_2_groupi_n_676 & csa_tree_add_69_2_groupi_n_654) | (csa_tree_add_69_2_groupi_n_654
    & csa_tree_add_69_2_groupi_n_932)));
 assign csa_tree_add_69_2_groupi_n_1121 = (csa_tree_add_69_2_groupi_n_676 ^ (csa_tree_add_69_2_groupi_n_654
    ^ csa_tree_add_69_2_groupi_n_932));
 assign csa_tree_add_69_2_groupi_n_1118 = ((csa_tree_add_69_2_groupi_n_856 & csa_tree_add_69_2_groupi_n_779)
    | ((csa_tree_add_69_2_groupi_n_779 & csa_tree_add_69_2_groupi_n_817) | (csa_tree_add_69_2_groupi_n_817
    & csa_tree_add_69_2_groupi_n_856)));
 assign csa_tree_add_69_2_groupi_n_1119 = (csa_tree_add_69_2_groupi_n_779 ^ (csa_tree_add_69_2_groupi_n_817
    ^ csa_tree_add_69_2_groupi_n_856));
 assign csa_tree_add_69_2_groupi_n_1116 = ((csa_tree_add_69_2_groupi_n_930 & csa_tree_add_69_2_groupi_n_669)
    | ((csa_tree_add_69_2_groupi_n_669 & csa_tree_add_69_2_groupi_n_657) | (csa_tree_add_69_2_groupi_n_657
    & csa_tree_add_69_2_groupi_n_930)));
 assign csa_tree_add_69_2_groupi_n_1117 = (csa_tree_add_69_2_groupi_n_669 ^ (csa_tree_add_69_2_groupi_n_657
    ^ csa_tree_add_69_2_groupi_n_930));
 assign csa_tree_add_69_2_groupi_n_1114 = ((csa_tree_add_69_2_groupi_n_706 & csa_tree_add_69_2_groupi_n_720)
    | ((csa_tree_add_69_2_groupi_n_720 & csa_tree_add_69_2_groupi_n_915) | (csa_tree_add_69_2_groupi_n_915
    & csa_tree_add_69_2_groupi_n_706)));
 assign csa_tree_add_69_2_groupi_n_1115 = (csa_tree_add_69_2_groupi_n_720 ^ (csa_tree_add_69_2_groupi_n_915
    ^ csa_tree_add_69_2_groupi_n_706));
 assign csa_tree_add_69_2_groupi_n_1112 = ((csa_tree_add_69_2_groupi_n_702 & csa_tree_add_69_2_groupi_n_724)
    | ((csa_tree_add_69_2_groupi_n_724 & csa_tree_add_69_2_groupi_n_885) | (csa_tree_add_69_2_groupi_n_885
    & csa_tree_add_69_2_groupi_n_702)));
 assign csa_tree_add_69_2_groupi_n_1113 = (csa_tree_add_69_2_groupi_n_724 ^ (csa_tree_add_69_2_groupi_n_885
    ^ csa_tree_add_69_2_groupi_n_702));
 assign csa_tree_add_69_2_groupi_n_1110 = ((csa_tree_add_69_2_groupi_n_927 & csa_tree_add_69_2_groupi_n_673)
    | ((csa_tree_add_69_2_groupi_n_673 & csa_tree_add_69_2_groupi_n_667) | (csa_tree_add_69_2_groupi_n_667
    & csa_tree_add_69_2_groupi_n_927)));
 assign csa_tree_add_69_2_groupi_n_1111 = (csa_tree_add_69_2_groupi_n_673 ^ (csa_tree_add_69_2_groupi_n_667
    ^ csa_tree_add_69_2_groupi_n_927));
 assign csa_tree_add_69_2_groupi_n_1108 = ((csa_tree_add_69_2_groupi_n_928 & csa_tree_add_69_2_groupi_n_718)
    | ((csa_tree_add_69_2_groupi_n_718 & csa_tree_add_69_2_groupi_n_671) | (csa_tree_add_69_2_groupi_n_671
    & csa_tree_add_69_2_groupi_n_928)));
 assign csa_tree_add_69_2_groupi_n_1109 = (csa_tree_add_69_2_groupi_n_718 ^ (csa_tree_add_69_2_groupi_n_671
    ^ csa_tree_add_69_2_groupi_n_928));
 assign csa_tree_add_69_2_groupi_n_1106 = ((csa_tree_add_69_2_groupi_n_852 & csa_tree_add_69_2_groupi_n_799)
    | ((csa_tree_add_69_2_groupi_n_799 & csa_tree_add_69_2_groupi_n_798) | (csa_tree_add_69_2_groupi_n_798
    & csa_tree_add_69_2_groupi_n_852)));
 assign csa_tree_add_69_2_groupi_n_1107 = (csa_tree_add_69_2_groupi_n_799 ^ (csa_tree_add_69_2_groupi_n_798
    ^ csa_tree_add_69_2_groupi_n_852));
 assign csa_tree_add_69_2_groupi_n_1104 = ((csa_tree_add_69_2_groupi_n_929 & csa_tree_add_69_2_groupi_n_659)
    | ((csa_tree_add_69_2_groupi_n_659 & csa_tree_add_69_2_groupi_n_660) | (csa_tree_add_69_2_groupi_n_660
    & csa_tree_add_69_2_groupi_n_929)));
 assign csa_tree_add_69_2_groupi_n_1105 = (csa_tree_add_69_2_groupi_n_659 ^ (csa_tree_add_69_2_groupi_n_660
    ^ csa_tree_add_69_2_groupi_n_929));
 assign csa_tree_add_69_2_groupi_n_1102 = ((csa_tree_add_69_2_groupi_n_840 & csa_tree_add_69_2_groupi_n_827)
    | ((csa_tree_add_69_2_groupi_n_827 & csa_tree_add_69_2_groupi_n_810) | (csa_tree_add_69_2_groupi_n_810
    & csa_tree_add_69_2_groupi_n_840)));
 assign csa_tree_add_69_2_groupi_n_1103 = (csa_tree_add_69_2_groupi_n_827 ^ (csa_tree_add_69_2_groupi_n_810
    ^ csa_tree_add_69_2_groupi_n_840));
 assign csa_tree_add_69_2_groupi_n_1100 = ((csa_tree_add_69_2_groupi_n_857 & csa_tree_add_69_2_groupi_n_773)
    | ((csa_tree_add_69_2_groupi_n_773 & csa_tree_add_69_2_groupi_n_818) | (csa_tree_add_69_2_groupi_n_818
    & csa_tree_add_69_2_groupi_n_857)));
 assign csa_tree_add_69_2_groupi_n_1101 = (csa_tree_add_69_2_groupi_n_773 ^ (csa_tree_add_69_2_groupi_n_818
    ^ csa_tree_add_69_2_groupi_n_857));
 assign csa_tree_add_69_2_groupi_n_1098 = ((csa_tree_add_69_2_groupi_n_842 & csa_tree_add_69_2_groupi_n_832)
    | ((csa_tree_add_69_2_groupi_n_832 & csa_tree_add_69_2_groupi_n_803) | (csa_tree_add_69_2_groupi_n_803
    & csa_tree_add_69_2_groupi_n_842)));
 assign csa_tree_add_69_2_groupi_n_1099 = (csa_tree_add_69_2_groupi_n_832 ^ (csa_tree_add_69_2_groupi_n_803
    ^ csa_tree_add_69_2_groupi_n_842));
 assign csa_tree_add_69_2_groupi_n_1097 = ~(csa_tree_add_69_2_groupi_n_1009 ^ csa_tree_add_69_2_groupi_n_1005);
 assign csa_tree_add_69_2_groupi_n_1096 = ~((csa_tree_add_69_2_groupi_n_1074 & ~csa_tree_add_69_2_groupi_n_1071)
    | (n_448 & csa_tree_add_69_2_groupi_n_1071));
 assign csa_tree_add_69_2_groupi_n_1142 = ~(csa_tree_add_69_2_groupi_n_998 | (csa_tree_add_69_2_groupi_n_983
    & csa_tree_add_69_2_groupi_n_997));
 assign csa_tree_add_69_2_groupi_n_1141 = ~(csa_tree_add_69_2_groupi_n_1081 | csa_tree_add_69_2_groupi_n_1000);
 assign csa_tree_add_69_2_groupi_n_1140 = ~(csa_tree_add_69_2_groupi_n_26 | csa_tree_add_69_2_groupi_n_23);
 assign csa_tree_add_69_2_groupi_n_1139 = ~((csa_tree_add_69_2_groupi_n_713 & ~csa_tree_add_69_2_groupi_n_1007)
    | (csa_tree_add_69_2_groupi_n_712 & csa_tree_add_69_2_groupi_n_1007));
 assign csa_tree_add_69_2_groupi_n_1138 = ~(csa_tree_add_69_2_groupi_n_1082 | csa_tree_add_69_2_groupi_n_32);
 assign csa_tree_add_69_2_groupi_n_1095 = ~(csa_tree_add_69_2_groupi_n_1008 ^ csa_tree_add_69_2_groupi_n_983);
 assign csa_tree_add_69_2_groupi_n_1094 = ~(csa_tree_add_69_2_groupi_n_1083 | ~csa_tree_add_69_2_groupi_n_964);
 assign csa_tree_add_69_2_groupi_n_1093 = ~(csa_tree_add_69_2_groupi_n_1079 | csa_tree_add_69_2_groupi_n_31);
 assign csa_tree_add_69_2_groupi_n_1092 = (csa_tree_add_69_2_groupi_n_1018 ^ csa_tree_add_69_2_groupi_n_875);
 assign csa_tree_add_69_2_groupi_n_1091 = ~(csa_tree_add_69_2_groupi_n_1017 ^ csa_tree_add_69_2_groupi_n_978);
 assign csa_tree_add_69_2_groupi_n_1089 = (csa_tree_add_69_2_groupi_n_1019 ^ csa_tree_add_69_2_groupi_n_977);
 assign csa_tree_add_69_2_groupi_n_1088 = ~(csa_tree_add_69_2_groupi_n_976 ^ (csa_tree_add_69_2_groupi_n_863
    ^ csa_tree_add_69_2_groupi_n_1072));
 assign csa_tree_add_69_2_groupi_n_1090 = ~(csa_tree_add_69_2_groupi_n_1078 | csa_tree_add_69_2_groupi_n_28);
 assign csa_tree_add_69_2_groupi_n_1087 = ~(csa_tree_add_69_2_groupi_n_991 & (csa_tree_add_69_2_groupi_n_990
    | csa_tree_add_69_2_groupi_n_979));
 assign csa_tree_add_69_2_groupi_n_1085 = ((csa_tree_add_69_2_groupi_n_858 & csa_tree_add_69_2_groupi_n_615)
    | ((csa_tree_add_69_2_groupi_n_615 & csa_tree_add_69_2_groupi_n_616) | (csa_tree_add_69_2_groupi_n_616
    & csa_tree_add_69_2_groupi_n_858)));
 assign csa_tree_add_69_2_groupi_n_1086 = (csa_tree_add_69_2_groupi_n_615 ^ (csa_tree_add_69_2_groupi_n_616
    ^ csa_tree_add_69_2_groupi_n_858));
 assign csa_tree_add_69_2_groupi_n_1084 = ~(csa_tree_add_69_2_groupi_n_1071 | ~n_448);
 assign csa_tree_add_69_2_groupi_n_1083 = ~(csa_tree_add_69_2_groupi_n_1012 | csa_tree_add_69_2_groupi_n_965);
 assign csa_tree_add_69_2_groupi_n_1082 = ~(csa_tree_add_69_2_groupi_n_989 | csa_tree_add_69_2_groupi_n_713);
 assign csa_tree_add_69_2_groupi_n_1081 = ~(csa_tree_add_69_2_groupi_n_1073 | (csa_tree_add_69_2_groupi_n_864
    & csa_tree_add_69_2_groupi_n_976));
 assign csa_tree_add_69_2_groupi_n_1079 = ~(csa_tree_add_69_2_groupi_n_993 | csa_tree_add_69_2_groupi_n_977);
 assign csa_tree_add_69_2_groupi_n_1078 = ~(csa_tree_add_69_2_groupi_n_988 | csa_tree_add_69_2_groupi_n_875);
 assign csa_tree_add_69_2_groupi_n_1077 = ~(csa_tree_add_69_2_groupi_n_1010 ^ csa_tree_add_69_2_groupi_n_960);
 assign csa_tree_add_69_2_groupi_n_1076 = ~(csa_tree_add_69_2_groupi_n_1016 ^ csa_tree_add_69_2_groupi_n_961);
 assign csa_tree_add_69_2_groupi_n_1075 = ~(csa_tree_add_69_2_groupi_n_1020 ^ csa_tree_add_69_2_groupi_n_867);
 assign csa_tree_add_69_2_groupi_n_1074 = ~n_448;
 assign csa_tree_add_69_2_groupi_n_1073 = ~csa_tree_add_69_2_groupi_n_1072;
 assign csa_tree_add_69_2_groupi_n_1069 = (csa_tree_add_69_2_groupi_n_954 & csa_tree_add_69_2_groupi_n_698);
 assign csa_tree_add_69_2_groupi_n_1070 = (csa_tree_add_69_2_groupi_n_954 ^ csa_tree_add_69_2_groupi_n_698);
 assign csa_tree_add_69_2_groupi_n_1067 = (csa_tree_add_69_2_groupi_n_935 & csa_tree_add_69_2_groupi_n_683);
 assign csa_tree_add_69_2_groupi_n_1068 = (csa_tree_add_69_2_groupi_n_935 ^ csa_tree_add_69_2_groupi_n_683);
 assign csa_tree_add_69_2_groupi_n_1065 = (csa_tree_add_69_2_groupi_n_936 & csa_tree_add_69_2_groupi_n_703);
 assign csa_tree_add_69_2_groupi_n_1066 = (csa_tree_add_69_2_groupi_n_936 ^ csa_tree_add_69_2_groupi_n_703);
 assign csa_tree_add_69_2_groupi_n_1063 = (csa_tree_add_69_2_groupi_n_947 & csa_tree_add_69_2_groupi_n_687);
 assign csa_tree_add_69_2_groupi_n_1064 = (csa_tree_add_69_2_groupi_n_947 ^ csa_tree_add_69_2_groupi_n_687);
 assign csa_tree_add_69_2_groupi_n_1061 = (csa_tree_add_69_2_groupi_n_938 & csa_tree_add_69_2_groupi_n_691);
 assign csa_tree_add_69_2_groupi_n_1062 = (csa_tree_add_69_2_groupi_n_938 ^ csa_tree_add_69_2_groupi_n_691);
 assign csa_tree_add_69_2_groupi_n_1059 = (csa_tree_add_69_2_groupi_n_953 & csa_tree_add_69_2_groupi_n_678);
 assign csa_tree_add_69_2_groupi_n_1060 = (csa_tree_add_69_2_groupi_n_953 ^ csa_tree_add_69_2_groupi_n_678);
 assign csa_tree_add_69_2_groupi_n_1057 = (csa_tree_add_69_2_groupi_n_701 & csa_tree_add_69_2_groupi_n_941);
 assign csa_tree_add_69_2_groupi_n_1058 = (csa_tree_add_69_2_groupi_n_701 ^ csa_tree_add_69_2_groupi_n_941);
 assign csa_tree_add_69_2_groupi_n_1055 = (csa_tree_add_69_2_groupi_n_926 & csa_tree_add_69_2_groupi_n_680);
 assign csa_tree_add_69_2_groupi_n_1056 = (csa_tree_add_69_2_groupi_n_926 ^ csa_tree_add_69_2_groupi_n_680);
 assign csa_tree_add_69_2_groupi_n_1053 = (csa_tree_add_69_2_groupi_n_952 & csa_tree_add_69_2_groupi_n_682);
 assign csa_tree_add_69_2_groupi_n_1054 = (csa_tree_add_69_2_groupi_n_952 ^ csa_tree_add_69_2_groupi_n_682);
 assign csa_tree_add_69_2_groupi_n_1051 = (csa_tree_add_69_2_groupi_n_957 & csa_tree_add_69_2_groupi_n_679);
 assign csa_tree_add_69_2_groupi_n_1052 = (csa_tree_add_69_2_groupi_n_957 ^ csa_tree_add_69_2_groupi_n_679);
 assign csa_tree_add_69_2_groupi_n_1049 = (csa_tree_add_69_2_groupi_n_931 & csa_tree_add_69_2_groupi_n_681);
 assign csa_tree_add_69_2_groupi_n_1050 = (csa_tree_add_69_2_groupi_n_931 ^ csa_tree_add_69_2_groupi_n_681);
 assign csa_tree_add_69_2_groupi_n_1047 = (csa_tree_add_69_2_groupi_n_937 & csa_tree_add_69_2_groupi_n_705);
 assign csa_tree_add_69_2_groupi_n_1048 = (csa_tree_add_69_2_groupi_n_937 ^ csa_tree_add_69_2_groupi_n_705);
 assign csa_tree_add_69_2_groupi_n_1045 = (csa_tree_add_69_2_groupi_n_951 & csa_tree_add_69_2_groupi_n_685);
 assign csa_tree_add_69_2_groupi_n_1046 = (csa_tree_add_69_2_groupi_n_951 ^ csa_tree_add_69_2_groupi_n_685);
 assign csa_tree_add_69_2_groupi_n_1043 = (csa_tree_add_69_2_groupi_n_949 & csa_tree_add_69_2_groupi_n_690);
 assign csa_tree_add_69_2_groupi_n_1044 = (csa_tree_add_69_2_groupi_n_949 ^ csa_tree_add_69_2_groupi_n_690);
 assign csa_tree_add_69_2_groupi_n_1041 = (csa_tree_add_69_2_groupi_n_944 & csa_tree_add_69_2_groupi_n_697);
 assign csa_tree_add_69_2_groupi_n_1042 = (csa_tree_add_69_2_groupi_n_944 ^ csa_tree_add_69_2_groupi_n_697);
 assign csa_tree_add_69_2_groupi_n_1039 = (csa_tree_add_69_2_groupi_n_940 & csa_tree_add_69_2_groupi_n_699);
 assign csa_tree_add_69_2_groupi_n_1040 = (csa_tree_add_69_2_groupi_n_940 ^ csa_tree_add_69_2_groupi_n_699);
 assign csa_tree_add_69_2_groupi_n_1037 = (csa_tree_add_69_2_groupi_n_950 & csa_tree_add_69_2_groupi_n_684);
 assign csa_tree_add_69_2_groupi_n_1038 = (csa_tree_add_69_2_groupi_n_950 ^ csa_tree_add_69_2_groupi_n_684);
 assign csa_tree_add_69_2_groupi_n_1072 = (csa_tree_add_69_2_groupi_n_946 & csa_tree_add_69_2_groupi_n_688);
 assign csa_tree_add_69_2_groupi_n_1036 = (csa_tree_add_69_2_groupi_n_946 ^ csa_tree_add_69_2_groupi_n_688);
 assign csa_tree_add_69_2_groupi_n_1071 = ((csa_tree_add_69_2_groupi_n_837 & csa_tree_add_69_2_groupi_n_558)
    | ((csa_tree_add_69_2_groupi_n_558 & csa_tree_add_69_2_groupi_n_559) | (csa_tree_add_69_2_groupi_n_559
    & csa_tree_add_69_2_groupi_n_837)));
 assign csa_tree_add_69_2_groupi_n_1035 = (csa_tree_add_69_2_groupi_n_558 ^ (csa_tree_add_69_2_groupi_n_559
    ^ csa_tree_add_69_2_groupi_n_837));
 assign csa_tree_add_69_2_groupi_n_1033 = (csa_tree_add_69_2_groupi_n_956 & csa_tree_add_69_2_groupi_n_692);
 assign csa_tree_add_69_2_groupi_n_1034 = (csa_tree_add_69_2_groupi_n_956 ^ csa_tree_add_69_2_groupi_n_692);
 assign csa_tree_add_69_2_groupi_n_1031 = (csa_tree_add_69_2_groupi_n_948 & csa_tree_add_69_2_groupi_n_686);
 assign csa_tree_add_69_2_groupi_n_1032 = (csa_tree_add_69_2_groupi_n_948 ^ csa_tree_add_69_2_groupi_n_686);
 assign csa_tree_add_69_2_groupi_n_1029 = (csa_tree_add_69_2_groupi_n_955 & csa_tree_add_69_2_groupi_n_677);
 assign csa_tree_add_69_2_groupi_n_1030 = (csa_tree_add_69_2_groupi_n_955 ^ csa_tree_add_69_2_groupi_n_677);
 assign csa_tree_add_69_2_groupi_n_1027 = (csa_tree_add_69_2_groupi_n_943 & csa_tree_add_69_2_groupi_n_696);
 assign csa_tree_add_69_2_groupi_n_1028 = (csa_tree_add_69_2_groupi_n_943 ^ csa_tree_add_69_2_groupi_n_696);
 assign csa_tree_add_69_2_groupi_n_1023 = ~(csa_tree_add_69_2_groupi_n_994 & ~csa_tree_add_69_2_groupi_n_862);
 assign csa_tree_add_69_2_groupi_n_1025 = ~(csa_tree_add_69_2_groupi_n_1021 | csa_tree_add_69_2_groupi_n_29);
 assign csa_tree_add_69_2_groupi_n_1024 = ~(csa_tree_add_69_2_groupi_n_1001 & (csa_tree_add_69_2_groupi_n_24
    | csa_tree_add_69_2_groupi_n_980));
 assign csa_tree_add_69_2_groupi_n_1021 = ~(csa_tree_add_69_2_groupi_n_992 | csa_tree_add_69_2_groupi_n_877);
 assign csa_tree_add_69_2_groupi_n_1020 = ~((csa_tree_add_69_2_groupi_n_876 & ~csa_tree_add_69_2_groupi_n_868)
    | (csa_tree_add_69_2_groupi_n_877 & csa_tree_add_69_2_groupi_n_868));
 assign csa_tree_add_69_2_groupi_n_1019 = ~((csa_tree_add_69_2_groupi_n_870 & ~csa_tree_add_69_2_groupi_n_968)
    | (csa_tree_add_69_2_groupi_n_869 & csa_tree_add_69_2_groupi_n_968));
 assign csa_tree_add_69_2_groupi_n_1018 = ~((csa_tree_add_69_2_groupi_n_860 & ~csa_tree_add_69_2_groupi_n_866)
    | (csa_tree_add_69_2_groupi_n_861 & csa_tree_add_69_2_groupi_n_866));
 assign csa_tree_add_69_2_groupi_n_1017 = ~((csa_tree_add_69_2_groupi_n_872 & ~csa_tree_add_69_2_groupi_n_873)
    | (csa_tree_add_69_2_groupi_n_871 & csa_tree_add_69_2_groupi_n_873));
 assign csa_tree_add_69_2_groupi_n_1016 = ~(csa_tree_add_69_2_groupi_n_962 ^ csa_tree_add_69_2_groupi_n_708);
 assign csa_tree_add_69_2_groupi_n_1015 = ~(csa_tree_add_69_2_groupi_n_1005 & (csa_tree_add_69_2_groupi_n_716
    | csa_tree_add_69_2_groupi_n_984));
 assign csa_tree_add_69_2_groupi_n_1010 = ~(csa_tree_add_69_2_groupi_n_730 ^ csa_tree_add_69_2_groupi_n_959);
 assign csa_tree_add_69_2_groupi_n_1009 = ~(csa_tree_add_69_2_groupi_n_963 ^ csa_tree_add_69_2_groupi_n_958);
 assign csa_tree_add_69_2_groupi_n_1013 = ~(csa_tree_add_69_2_groupi_n_999 | (csa_tree_add_69_2_groupi_n_711
    & csa_tree_add_69_2_groupi_n_980));
 assign csa_tree_add_69_2_groupi_n_1008 = ~((csa_tree_add_69_2_groupi_n_974 & ~csa_tree_add_69_2_groupi_n_972)
    | (csa_tree_add_69_2_groupi_n_973 & csa_tree_add_69_2_groupi_n_972));
 assign csa_tree_add_69_2_groupi_n_1007 = ~((csa_tree_add_69_2_groupi_n_970 & ~csa_tree_add_69_2_groupi_n_969)
    | (csa_tree_add_69_2_groupi_n_971 & csa_tree_add_69_2_groupi_n_969));
 assign csa_tree_add_69_2_groupi_n_1012 = ~(csa_tree_add_69_2_groupi_n_981 ^ csa_tree_add_69_2_groupi_n_581);
 assign csa_tree_add_69_2_groupi_n_1011 = ~(csa_tree_add_69_2_groupi_n_987 & ~(csa_tree_add_69_2_groupi_n_431
    & csa_tree_add_69_2_groupi_n_430));
 assign csa_tree_add_69_2_groupi_n_1003 = (csa_tree_add_69_2_groupi_n_617 & csa_tree_add_69_2_groupi_n_619);
 assign csa_tree_add_69_2_groupi_n_1004 = (csa_tree_add_69_2_groupi_n_617 ^ csa_tree_add_69_2_groupi_n_619);
 assign csa_tree_add_69_2_groupi_n_1001 = ~(csa_tree_add_69_2_groupi_n_711 & csa_tree_add_69_2_groupi_n_967);
 assign csa_tree_add_69_2_groupi_n_1000 = ~(csa_tree_add_69_2_groupi_n_976 | ~csa_tree_add_69_2_groupi_n_863);
 assign csa_tree_add_69_2_groupi_n_999 = ~(csa_tree_add_69_2_groupi_n_771 | (csa_tree_add_69_2_groupi_n_77
    | csa_tree_add_69_2_groupi_n_711));
 assign csa_tree_add_69_2_groupi_n_998 = ~(csa_tree_add_69_2_groupi_n_974 | csa_tree_add_69_2_groupi_n_972);
 assign csa_tree_add_69_2_groupi_n_997 = ~(csa_tree_add_69_2_groupi_n_974 & csa_tree_add_69_2_groupi_n_972);
 assign csa_tree_add_69_2_groupi_n_1005 = ~(csa_tree_add_69_2_groupi_n_716 & csa_tree_add_69_2_groupi_n_984);
 assign csa_tree_add_69_2_groupi_n_995 = ~(csa_tree_add_69_2_groupi_n_982 & csa_tree_add_69_2_groupi_n_714);
 assign csa_tree_add_69_2_groupi_n_993 = ~(csa_tree_add_69_2_groupi_n_968 | csa_tree_add_69_2_groupi_n_870);
 assign csa_tree_add_69_2_groupi_n_992 = ~(csa_tree_add_69_2_groupi_n_867 | csa_tree_add_69_2_groupi_n_868);
 assign csa_tree_add_69_2_groupi_n_991 = ~(csa_tree_add_69_2_groupi_n_874 & csa_tree_add_69_2_groupi_n_872);
 assign csa_tree_add_69_2_groupi_n_990 = ~(csa_tree_add_69_2_groupi_n_874 | csa_tree_add_69_2_groupi_n_872);
 assign csa_tree_add_69_2_groupi_n_989 = ~(csa_tree_add_69_2_groupi_n_969 | csa_tree_add_69_2_groupi_n_971);
 assign csa_tree_add_69_2_groupi_n_988 = ~(csa_tree_add_69_2_groupi_n_866 | ~csa_tree_add_69_2_groupi_n_861);
 assign csa_tree_add_69_2_groupi_n_987 = ~(csa_tree_add_69_2_groupi_n_981 & csa_tree_add_69_2_groupi_n_561);
 assign csa_tree_add_69_2_groupi_n_994 = (csa_tree_add_69_2_groupi_n_618 ^ csa_tree_add_69_2_groupi_n_715);
 assign csa_tree_add_69_2_groupi_n_985 = ~(csa_tree_add_69_2_groupi_n_878 | csa_tree_add_69_2_groupi_n_880);
 assign csa_tree_add_69_2_groupi_n_979 = ~csa_tree_add_69_2_groupi_n_978;
 assign csa_tree_add_69_2_groupi_n_974 = ~csa_tree_add_69_2_groupi_n_973;
 assign csa_tree_add_69_2_groupi_n_970 = ~csa_tree_add_69_2_groupi_n_971;
 assign csa_tree_add_69_2_groupi_n_967 = ~csa_tree_add_69_2_groupi_n_966;
 assign csa_tree_add_69_2_groupi_n_965 = ~(csa_tree_add_69_2_groupi_n_709 | csa_tree_add_69_2_groupi_n_653);
 assign csa_tree_add_69_2_groupi_n_964 = ~(csa_tree_add_69_2_groupi_n_709 & csa_tree_add_69_2_groupi_n_653);
 assign csa_tree_add_69_2_groupi_n_963 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_531)
    & (n_487 | csa_tree_add_69_2_groupi_n_421));
 assign csa_tree_add_69_2_groupi_n_962 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_541)
    & (n_488 | csa_tree_add_69_2_groupi_n_422));
 assign csa_tree_add_69_2_groupi_n_961 = ~((n_456 | csa_tree_add_69_2_groupi_n_538) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_134));
 assign csa_tree_add_69_2_groupi_n_960 = ~((csa_tree_add_69_2_groupi_n_652 & csa_tree_add_69_2_groupi_n_506)
    | (n_485 & csa_tree_add_69_2_groupi_n_414));
 assign csa_tree_add_69_2_groupi_n_959 = ~((csa_tree_add_69_2_groupi_n_650 & csa_tree_add_69_2_groupi_n_504)
    | (n_486 & csa_tree_add_69_2_groupi_n_415));
 assign csa_tree_add_69_2_groupi_n_984 = ~(csa_tree_add_69_2_groupi_n_227 & ~(csa_tree_add_69_2_groupi_n_642
    & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_958 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_529)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_420));
 assign csa_tree_add_69_2_groupi_n_957 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_439)
    & (csa_tree_add_69_2_groupi_n_524 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_983 = ~(csa_tree_add_69_2_groupi_n_766 & csa_tree_add_69_2_groupi_n_562);
 assign csa_tree_add_69_2_groupi_n_956 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_450)
    & (csa_tree_add_69_2_groupi_n_439 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_955 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_447)
    & (csa_tree_add_69_2_groupi_n_459 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_954 = ~(csa_tree_add_69_2_groupi_n_554 & ~(csa_tree_add_69_2_groupi_n_642
    & csa_tree_add_69_2_groupi_n_441));
 assign csa_tree_add_69_2_groupi_n_953 = ~(csa_tree_add_69_2_groupi_n_570 & ~(csa_tree_add_69_2_groupi_n_642
    & csa_tree_add_69_2_groupi_n_446));
 assign csa_tree_add_69_2_groupi_n_952 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_302)
    & (csa_tree_add_69_2_groupi_n_447 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_951 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_498)
    & (csa_tree_add_69_2_groupi_n_516 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_950 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_516)
    & (csa_tree_add_69_2_groupi_n_515 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_949 = ~(csa_tree_add_69_2_groupi_n_551 & ~(csa_tree_add_69_2_groupi_n_642
    & n_483));
 assign csa_tree_add_69_2_groupi_n_948 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_468)
    & (csa_tree_add_69_2_groupi_n_437 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_982 = ~(csa_tree_add_69_2_groupi_n_743 & csa_tree_add_69_2_groupi_n_571);
 assign csa_tree_add_69_2_groupi_n_947 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_436)
    & (csa_tree_add_69_2_groupi_n_302 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_946 = ~(csa_tree_add_69_2_groupi_n_767 & csa_tree_add_69_2_groupi_n_556);
 assign csa_tree_add_69_2_groupi_n_945 = ~(csa_tree_add_69_2_groupi_n_772 & ~csa_tree_add_69_2_groupi_n_99);
 assign csa_tree_add_69_2_groupi_n_944 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_460)
    & (csa_tree_add_69_2_groupi_n_436 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_981 = ~(csa_tree_add_69_2_groupi_n_764 & csa_tree_add_69_2_groupi_n_553);
 assign csa_tree_add_69_2_groupi_n_943 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_452)
    & (csa_tree_add_69_2_groupi_n_303 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_980 = ~(csa_tree_add_69_2_groupi_n_770 & n_382);
 assign csa_tree_add_69_2_groupi_n_942 = ~(n_487 | (csa_tree_add_69_2_groupi_n_100 | csa_tree_add_69_2_groupi_n_715));
 assign csa_tree_add_69_2_groupi_n_941 = ~(csa_tree_add_69_2_groupi_n_227 & (csa_tree_add_69_2_groupi_n_641
    | csa_tree_add_69_2_groupi_n_526));
 assign csa_tree_add_69_2_groupi_n_940 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_515)
    & (csa_tree_add_69_2_groupi_n_502 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_939 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_510)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_529));
 assign csa_tree_add_69_2_groupi_n_938 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_437)
    & (csa_tree_add_69_2_groupi_n_498 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_937 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_502)
    & (csa_tree_add_69_2_groupi_n_525 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_936 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_525)
    & (csa_tree_add_69_2_groupi_n_526 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_935 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_303)
    & (csa_tree_add_69_2_groupi_n_460 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_934 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_334)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_313));
 assign csa_tree_add_69_2_groupi_n_933 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_319)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_309));
 assign csa_tree_add_69_2_groupi_n_932 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_316)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_348));
 assign csa_tree_add_69_2_groupi_n_931 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_524)
    & (csa_tree_add_69_2_groupi_n_452 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_930 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_331)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_344));
 assign csa_tree_add_69_2_groupi_n_978 = ~(csa_tree_add_69_2_groupi_n_639 & ~(csa_tree_add_69_2_groupi_n_650
    & n_508));
 assign csa_tree_add_69_2_groupi_n_929 = ~(csa_tree_add_69_2_groupi_n_761 & csa_tree_add_69_2_groupi_n_603);
 assign csa_tree_add_69_2_groupi_n_977 = ~(csa_tree_add_69_2_groupi_n_763 | csa_tree_add_69_2_groupi_n_12);
 assign csa_tree_add_69_2_groupi_n_928 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_306)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_339));
 assign csa_tree_add_69_2_groupi_n_927 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_309)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_340));
 assign csa_tree_add_69_2_groupi_n_926 = ~((csa_tree_add_69_2_groupi_n_641 | csa_tree_add_69_2_groupi_n_459)
    & (csa_tree_add_69_2_groupi_n_468 | csa_tree_add_69_2_groupi_n_71));
 assign csa_tree_add_69_2_groupi_n_925 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_513)
    & (n_488 | csa_tree_add_69_2_groupi_n_540));
 assign csa_tree_add_69_2_groupi_n_924 = ~(csa_tree_add_69_2_groupi_n_560 | (csa_tree_add_69_2_groupi_n_642
    & n_476));
 assign csa_tree_add_69_2_groupi_n_923 = ~(csa_tree_add_69_2_groupi_n_765 & csa_tree_add_69_2_groupi_n_563);
 assign csa_tree_add_69_2_groupi_n_976 = ~(csa_tree_add_69_2_groupi_n_735 & csa_tree_add_69_2_groupi_n_69);
 assign csa_tree_add_69_2_groupi_n_922 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_493)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_503));
 assign csa_tree_add_69_2_groupi_n_921 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_308)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_341));
 assign csa_tree_add_69_2_groupi_n_920 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_343)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_345));
 assign csa_tree_add_69_2_groupi_n_975 = ~(csa_tree_add_69_2_groupi_n_768 | csa_tree_add_69_2_groupi_n_555);
 assign csa_tree_add_69_2_groupi_n_919 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_347)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_308));
 assign csa_tree_add_69_2_groupi_n_918 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_337)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_323));
 assign csa_tree_add_69_2_groupi_n_917 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_349)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_321));
 assign csa_tree_add_69_2_groupi_n_916 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_348)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_334));
 assign csa_tree_add_69_2_groupi_n_915 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_344)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_350));
 assign csa_tree_add_69_2_groupi_n_973 = ~(csa_tree_add_69_2_groupi_n_733 | csa_tree_add_69_2_groupi_n_134);
 assign csa_tree_add_69_2_groupi_n_914 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_328)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_347));
 assign csa_tree_add_69_2_groupi_n_913 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_317)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_319));
 assign csa_tree_add_69_2_groupi_n_912 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_312)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_343));
 assign csa_tree_add_69_2_groupi_n_911 = ~((n_456 | csa_tree_add_69_2_groupi_n_537) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_536));
 assign csa_tree_add_69_2_groupi_n_910 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_330)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_328));
 assign csa_tree_add_69_2_groupi_n_909 = ~((n_456 | csa_tree_add_69_2_groupi_n_536) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_538));
 assign csa_tree_add_69_2_groupi_n_908 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_326)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_316));
 assign csa_tree_add_69_2_groupi_n_907 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_318)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_337));
 assign csa_tree_add_69_2_groupi_n_906 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_540)
    & (n_488 | csa_tree_add_69_2_groupi_n_530));
 assign csa_tree_add_69_2_groupi_n_905 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_333)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_330));
 assign csa_tree_add_69_2_groupi_n_904 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_340)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_493));
 assign csa_tree_add_69_2_groupi_n_903 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_345)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_310));
 assign csa_tree_add_69_2_groupi_n_902 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_305)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_312));
 assign csa_tree_add_69_2_groupi_n_901 = ~(csa_tree_add_69_2_groupi_n_762 & ~(n_486 & csa_tree_add_69_2_groupi_n_325));
 assign csa_tree_add_69_2_groupi_n_900 = ~(csa_tree_add_69_2_groupi_n_605 & ~(csa_tree_add_69_2_groupi_n_652
    & csa_tree_add_69_2_groupi_n_322));
 assign csa_tree_add_69_2_groupi_n_899 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_313)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_306));
 assign csa_tree_add_69_2_groupi_n_898 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_530)
    & (n_488 | csa_tree_add_69_2_groupi_n_541));
 assign csa_tree_add_69_2_groupi_n_972 = ~(csa_tree_add_69_2_groupi_n_732 & csa_tree_add_69_2_groupi_n_94);
 assign csa_tree_add_69_2_groupi_n_897 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_335)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_331));
 assign csa_tree_add_69_2_groupi_n_971 = ~(csa_tree_add_69_2_groupi_n_760 & csa_tree_add_69_2_groupi_n_635);
 assign csa_tree_add_69_2_groupi_n_969 = ~(csa_tree_add_69_2_groupi_n_759 & csa_tree_add_69_2_groupi_n_602);
 assign csa_tree_add_69_2_groupi_n_896 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_315)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_317));
 assign csa_tree_add_69_2_groupi_n_895 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_321)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_305));
 assign csa_tree_add_69_2_groupi_n_894 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_323)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_329));
 assign csa_tree_add_69_2_groupi_n_893 = ~(csa_tree_add_69_2_groupi_n_552 & ~(csa_tree_add_69_2_groupi_n_642
    & csa_tree_add_69_2_groupi_n_435));
 assign csa_tree_add_69_2_groupi_n_892 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_310)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_318));
 assign csa_tree_add_69_2_groupi_n_891 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_324)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_335));
 assign csa_tree_add_69_2_groupi_n_968 = ~(csa_tree_add_69_2_groupi_n_758 & csa_tree_add_69_2_groupi_n_611);
 assign csa_tree_add_69_2_groupi_n_890 = ~(csa_tree_add_69_2_groupi_n_757 & ~csa_tree_add_69_2_groupi_n_597);
 assign csa_tree_add_69_2_groupi_n_889 = ~(csa_tree_add_69_2_groupi_n_756 & csa_tree_add_69_2_groupi_n_598);
 assign csa_tree_add_69_2_groupi_n_888 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_329)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_494));
 assign csa_tree_add_69_2_groupi_n_887 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_494)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_505));
 assign csa_tree_add_69_2_groupi_n_886 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_339)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_324));
 assign csa_tree_add_69_2_groupi_n_885 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_350)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_346));
 assign csa_tree_add_69_2_groupi_n_884 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_509)
    & (n_487 | csa_tree_add_69_2_groupi_n_531));
 assign csa_tree_add_69_2_groupi_n_883 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_341)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_307));
 assign csa_tree_add_69_2_groupi_n_882 = ~((csa_tree_add_69_2_groupi_n_651 | csa_tree_add_69_2_groupi_n_307)
    & (csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_349));
 assign csa_tree_add_69_2_groupi_n_966 = ~(csa_tree_add_69_2_groupi_n_734 & csa_tree_add_69_2_groupi_n_67);
 assign csa_tree_add_69_2_groupi_n_881 = ~((n_456 | csa_tree_add_69_2_groupi_n_511) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_537));
 assign csa_tree_add_69_2_groupi_n_880 = ~csa_tree_add_69_2_groupi_n_879;
 assign csa_tree_add_69_2_groupi_n_877 = ~csa_tree_add_69_2_groupi_n_876;
 assign csa_tree_add_69_2_groupi_n_874 = ~csa_tree_add_69_2_groupi_n_873;
 assign csa_tree_add_69_2_groupi_n_872 = ~csa_tree_add_69_2_groupi_n_871;
 assign csa_tree_add_69_2_groupi_n_869 = ~csa_tree_add_69_2_groupi_n_870;
 assign csa_tree_add_69_2_groupi_n_864 = ~csa_tree_add_69_2_groupi_n_863;
 assign csa_tree_add_69_2_groupi_n_860 = ~csa_tree_add_69_2_groupi_n_861;
 assign csa_tree_add_69_2_groupi_n_859 = ~((csa_tree_add_69_2_groupi_n_649 | csa_tree_add_69_2_groupi_n_346)
    & (csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_315));
 assign csa_tree_add_69_2_groupi_n_858 = ~(csa_tree_add_69_2_groupi_n_737 & csa_tree_add_69_2_groupi_n_631);
 assign csa_tree_add_69_2_groupi_n_857 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_391)
    & (n_487 | csa_tree_add_69_2_groupi_n_373));
 assign csa_tree_add_69_2_groupi_n_879 = ~(csa_tree_add_69_2_groupi_n_738 & csa_tree_add_69_2_groupi_n_630);
 assign csa_tree_add_69_2_groupi_n_856 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_371)
    & (n_487 | csa_tree_add_69_2_groupi_n_393));
 assign csa_tree_add_69_2_groupi_n_855 = ~(csa_tree_add_69_2_groupi_n_740 | csa_tree_add_69_2_groupi_n_590);
 assign csa_tree_add_69_2_groupi_n_854 = ~(csa_tree_add_69_2_groupi_n_741 & csa_tree_add_69_2_groupi_n_18);
 assign csa_tree_add_69_2_groupi_n_878 = ~(csa_tree_add_69_2_groupi_n_769 | csa_tree_add_69_2_groupi_n_19);
 assign csa_tree_add_69_2_groupi_n_876 = ~(csa_tree_add_69_2_groupi_n_11 & csa_tree_add_69_2_groupi_n_604);
 assign csa_tree_add_69_2_groupi_n_853 = ~(csa_tree_add_69_2_groupi_n_594 & ~(csa_tree_add_69_2_groupi_n_92
    & n_491));
 assign csa_tree_add_69_2_groupi_n_852 = ~((n_456 | csa_tree_add_69_2_groupi_n_412) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_301));
 assign csa_tree_add_69_2_groupi_n_851 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_383)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_388));
 assign csa_tree_add_69_2_groupi_n_850 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_380)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_356));
 assign csa_tree_add_69_2_groupi_n_849 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_354)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_304));
 assign csa_tree_add_69_2_groupi_n_848 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_368)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_354));
 assign csa_tree_add_69_2_groupi_n_847 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_377)
    & (n_487 | csa_tree_add_69_2_groupi_n_371));
 assign csa_tree_add_69_2_groupi_n_846 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_507)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_510));
 assign csa_tree_add_69_2_groupi_n_845 = ~(csa_tree_add_69_2_groupi_n_753 & csa_tree_add_69_2_groupi_n_586);
 assign csa_tree_add_69_2_groupi_n_844 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_364)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_359));
 assign csa_tree_add_69_2_groupi_n_843 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_396)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_368));
 assign csa_tree_add_69_2_groupi_n_842 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_362)
    & (n_487 | csa_tree_add_69_2_groupi_n_363));
 assign csa_tree_add_69_2_groupi_n_841 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_496)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_507));
 assign csa_tree_add_69_2_groupi_n_840 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_363)
    & (n_487 | csa_tree_add_69_2_groupi_n_370));
 assign csa_tree_add_69_2_groupi_n_875 = ~(csa_tree_add_69_2_groupi_n_755 | csa_tree_add_69_2_groupi_n_596);
 assign csa_tree_add_69_2_groupi_n_839 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_359)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_496));
 assign csa_tree_add_69_2_groupi_n_838 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_372)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_369));
 assign csa_tree_add_69_2_groupi_n_837 = ~(csa_tree_add_69_2_groupi_n_748 & csa_tree_add_69_2_groupi_n_612);
 assign csa_tree_add_69_2_groupi_n_836 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_304)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_372));
 assign csa_tree_add_69_2_groupi_n_835 = ~(csa_tree_add_69_2_groupi_n_14 | csa_tree_add_69_2_groupi_n_591);
 assign csa_tree_add_69_2_groupi_n_834 = ~(csa_tree_add_69_2_groupi_n_595 | ~(csa_tree_add_69_2_groupi_n_647
    | csa_tree_add_69_2_groupi_n_390));
 assign csa_tree_add_69_2_groupi_n_833 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_357)
    & (n_487 | csa_tree_add_69_2_groupi_n_366));
 assign csa_tree_add_69_2_groupi_n_873 = ~(csa_tree_add_69_2_groupi_n_749 | csa_tree_add_69_2_groupi_n_607);
 assign csa_tree_add_69_2_groupi_n_832 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_356)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_355));
 assign csa_tree_add_69_2_groupi_n_871 = ~(csa_tree_add_69_2_groupi_n_15 | csa_tree_add_69_2_groupi_n_609);
 assign csa_tree_add_69_2_groupi_n_831 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_379)
    & (n_487 | csa_tree_add_69_2_groupi_n_357));
 assign csa_tree_add_69_2_groupi_n_830 = ~(csa_tree_add_69_2_groupi_n_746 & ~csa_tree_add_69_2_groupi_n_589);
 assign csa_tree_add_69_2_groupi_n_870 = ~(csa_tree_add_69_2_groupi_n_747 & csa_tree_add_69_2_groupi_n_599);
 assign csa_tree_add_69_2_groupi_n_868 = ~(n_452 & csa_tree_add_69_2_groupi_n_613);
 assign csa_tree_add_69_2_groupi_n_829 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_366)
    & (n_487 | csa_tree_add_69_2_groupi_n_377));
 assign csa_tree_add_69_2_groupi_n_867 = ~(csa_tree_add_69_2_groupi_n_750 & csa_tree_add_69_2_groupi_n_601);
 assign csa_tree_add_69_2_groupi_n_866 = ~(csa_tree_add_69_2_groupi_n_16 & csa_tree_add_69_2_groupi_n_600);
 assign csa_tree_add_69_2_groupi_n_828 = ~(csa_tree_add_69_2_groupi_n_745 & csa_tree_add_69_2_groupi_n_592);
 assign csa_tree_add_69_2_groupi_n_827 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_355)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_364));
 assign csa_tree_add_69_2_groupi_n_826 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_378)
    & (n_487 | csa_tree_add_69_2_groupi_n_495));
 assign csa_tree_add_69_2_groupi_n_825 = ~(csa_tree_add_69_2_groupi_n_754 & csa_tree_add_69_2_groupi_n_610);
 assign csa_tree_add_69_2_groupi_n_824 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_508)
    & (n_487 | csa_tree_add_69_2_groupi_n_509));
 assign csa_tree_add_69_2_groupi_n_823 = ~(csa_tree_add_69_2_groupi_n_13 & csa_tree_add_69_2_groupi_n_588);
 assign csa_tree_add_69_2_groupi_n_822 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_373)
    & (n_487 | csa_tree_add_69_2_groupi_n_392));
 assign csa_tree_add_69_2_groupi_n_821 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_369)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_376));
 assign csa_tree_add_69_2_groupi_n_820 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_392)
    & (n_487 | csa_tree_add_69_2_groupi_n_379));
 assign csa_tree_add_69_2_groupi_n_819 = ~((n_456 | csa_tree_add_69_2_groupi_n_410) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_295));
 assign csa_tree_add_69_2_groupi_n_818 = ~((n_456 | csa_tree_add_69_2_groupi_n_301) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_410));
 assign csa_tree_add_69_2_groupi_n_817 = ~((n_456 | csa_tree_add_69_2_groupi_n_401) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_398));
 assign csa_tree_add_69_2_groupi_n_816 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_370)
    & (n_487 | csa_tree_add_69_2_groupi_n_378));
 assign csa_tree_add_69_2_groupi_n_815 = ~((n_456 | csa_tree_add_69_2_groupi_n_300) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_412));
 assign csa_tree_add_69_2_groupi_n_814 = ~((n_456 | csa_tree_add_69_2_groupi_n_400) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_401));
 assign csa_tree_add_69_2_groupi_n_813 = ~((n_456 | csa_tree_add_69_2_groupi_n_497) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_512));
 assign csa_tree_add_69_2_groupi_n_812 = ~((n_456 | csa_tree_add_69_2_groupi_n_408) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_300));
 assign csa_tree_add_69_2_groupi_n_811 = ~(csa_tree_add_69_2_groupi_n_744 & csa_tree_add_69_2_groupi_n_606);
 assign csa_tree_add_69_2_groupi_n_810 = ~((n_456 | csa_tree_add_69_2_groupi_n_404) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_497));
 assign csa_tree_add_69_2_groupi_n_809 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_385)
    & (n_487 | csa_tree_add_69_2_groupi_n_387));
 assign csa_tree_add_69_2_groupi_n_808 = ~((n_456 | csa_tree_add_69_2_groupi_n_296) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_400));
 assign csa_tree_add_69_2_groupi_n_865 = ~(csa_tree_add_69_2_groupi_n_752 & csa_tree_add_69_2_groupi_n_17);
 assign csa_tree_add_69_2_groupi_n_807 = ~(csa_tree_add_69_2_groupi_n_608 & ~(csa_tree_add_69_2_groupi_n_92
    & n_492));
 assign csa_tree_add_69_2_groupi_n_806 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_393)
    & (n_487 | csa_tree_add_69_2_groupi_n_362));
 assign csa_tree_add_69_2_groupi_n_805 = ~((n_456 | csa_tree_add_69_2_groupi_n_512) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_511));
 assign csa_tree_add_69_2_groupi_n_804 = ~(csa_tree_add_69_2_groupi_n_587 & ~(csa_tree_add_69_2_groupi_n_92
    & n_494));
 assign csa_tree_add_69_2_groupi_n_803 = ~((n_456 | csa_tree_add_69_2_groupi_n_405) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_404));
 assign csa_tree_add_69_2_groupi_n_863 = ~(csa_tree_add_69_2_groupi_n_742 & csa_tree_add_69_2_groupi_n_593);
 assign csa_tree_add_69_2_groupi_n_802 = ~((n_456 | csa_tree_add_69_2_groupi_n_409) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_297));
 assign csa_tree_add_69_2_groupi_n_801 = ~((n_456 | csa_tree_add_69_2_groupi_n_297) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_296));
 assign csa_tree_add_69_2_groupi_n_800 = ~((n_456 | csa_tree_add_69_2_groupi_n_295) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_409));
 assign csa_tree_add_69_2_groupi_n_799 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_387)
    & (n_487 | csa_tree_add_69_2_groupi_n_391));
 assign csa_tree_add_69_2_groupi_n_798 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_388)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_394));
 assign csa_tree_add_69_2_groupi_n_797 = ~((n_456 | csa_tree_add_69_2_groupi_n_398) & (csa_tree_add_69_2_groupi_n_90
    | csa_tree_add_69_2_groupi_n_405));
 assign csa_tree_add_69_2_groupi_n_796 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_458)
    & (n_488 | csa_tree_add_69_2_groupi_n_527));
 assign csa_tree_add_69_2_groupi_n_795 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_465)
    & (n_488 | csa_tree_add_69_2_groupi_n_458));
 assign csa_tree_add_69_2_groupi_n_794 = ~(csa_tree_add_69_2_groupi_n_627 & ~(csa_tree_add_69_2_groupi_n_644
    & csa_tree_add_69_2_groupi_n_292));
 assign csa_tree_add_69_2_groupi_n_793 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_445)
    & (n_488 | csa_tree_add_69_2_groupi_n_358));
 assign csa_tree_add_69_2_groupi_n_792 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_461)
    & (n_488 | csa_tree_add_69_2_groupi_n_465));
 assign csa_tree_add_69_2_groupi_n_791 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_519)
    & (n_488 | csa_tree_add_69_2_groupi_n_451));
 assign csa_tree_add_69_2_groupi_n_790 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_462)
    & (n_488 | csa_tree_add_69_2_groupi_n_461));
 assign csa_tree_add_69_2_groupi_n_789 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_455)
    & (n_488 | csa_tree_add_69_2_groupi_n_445));
 assign csa_tree_add_69_2_groupi_n_788 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_454)
    & (n_488 | csa_tree_add_69_2_groupi_n_462));
 assign csa_tree_add_69_2_groupi_n_787 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_466)
    & (n_488 | csa_tree_add_69_2_groupi_n_443));
 assign csa_tree_add_69_2_groupi_n_786 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_499)
    & (n_488 | csa_tree_add_69_2_groupi_n_514));
 assign csa_tree_add_69_2_groupi_n_862 = ~(csa_tree_add_69_2_groupi_n_736 & csa_tree_add_69_2_groupi_n_626);
 assign csa_tree_add_69_2_groupi_n_785 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_451)
    & (n_488 | csa_tree_add_69_2_groupi_n_499));
 assign csa_tree_add_69_2_groupi_n_784 = ~(csa_tree_add_69_2_groupi_n_628 & ~(csa_tree_add_69_2_groupi_n_644
    & n_482));
 assign csa_tree_add_69_2_groupi_n_783 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_443)
    & (n_488 | csa_tree_add_69_2_groupi_n_455));
 assign csa_tree_add_69_2_groupi_n_782 = ~((csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_495)
    & (n_487 | csa_tree_add_69_2_groupi_n_508));
 assign csa_tree_add_69_2_groupi_n_781 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_514)
    & (n_488 | csa_tree_add_69_2_groupi_n_513));
 assign csa_tree_add_69_2_groupi_n_861 = ~(csa_tree_add_69_2_groupi_n_22 | csa_tree_add_69_2_groupi_n_20);
 assign csa_tree_add_69_2_groupi_n_780 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_522)
    & (n_488 | csa_tree_add_69_2_groupi_n_466));
 assign csa_tree_add_69_2_groupi_n_779 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_376)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_380));
 assign csa_tree_add_69_2_groupi_n_778 = ~(csa_tree_add_69_2_groupi_n_632 & ~(csa_tree_add_69_2_groupi_n_644
    & n_477));
 assign csa_tree_add_69_2_groupi_n_777 = ~(csa_tree_add_69_2_groupi_n_739 & csa_tree_add_69_2_groupi_n_633);
 assign csa_tree_add_69_2_groupi_n_776 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_527)
    & (n_488 | csa_tree_add_69_2_groupi_n_522));
 assign csa_tree_add_69_2_groupi_n_775 = ~(csa_tree_add_69_2_groupi_n_629 & ~(csa_tree_add_69_2_groupi_n_644
    & n_481));
 assign csa_tree_add_69_2_groupi_n_774 = ~((csa_tree_add_69_2_groupi_n_643 | csa_tree_add_69_2_groupi_n_358)
    & (n_488 | csa_tree_add_69_2_groupi_n_519));
 assign csa_tree_add_69_2_groupi_n_773 = ~((csa_tree_add_69_2_groupi_n_647 | csa_tree_add_69_2_groupi_n_394)
    & (csa_tree_add_69_2_groupi_n_577 | csa_tree_add_69_2_groupi_n_396));
 assign csa_tree_add_69_2_groupi_n_771 = ~csa_tree_add_69_2_groupi_n_770;
 assign csa_tree_add_69_2_groupi_n_769 = (csa_tree_add_69_2_groupi_n_92 & n_513);
 assign csa_tree_add_69_2_groupi_n_768 = (csa_tree_add_69_2_groupi_n_642 & n_462);
 assign csa_tree_add_69_2_groupi_n_767 = ~(csa_tree_add_69_2_groupi_n_642 & csa_tree_add_69_2_groupi_n_440);
 assign csa_tree_add_69_2_groupi_n_766 = ~(csa_tree_add_69_2_groupi_n_642 & n_460);
 assign csa_tree_add_69_2_groupi_n_765 = ~(csa_tree_add_69_2_groupi_n_642 & n_461);
 assign csa_tree_add_69_2_groupi_n_764 = ~(csa_tree_add_69_2_groupi_n_642 & n_489);
 assign csa_tree_add_69_2_groupi_n_763 = ~(csa_tree_add_69_2_groupi_n_651 | n_509);
 assign csa_tree_add_69_2_groupi_n_762 = ~(csa_tree_add_69_2_groupi_n_650 & n_510);
 assign csa_tree_add_69_2_groupi_n_761 = ~(csa_tree_add_69_2_groupi_n_652 & n_505);
 assign csa_tree_add_69_2_groupi_n_760 = ~(csa_tree_add_69_2_groupi_n_652 & n_511);
 assign csa_tree_add_69_2_groupi_n_759 = ~(csa_tree_add_69_2_groupi_n_650 & n_504);
 assign csa_tree_add_69_2_groupi_n_758 = ~(csa_tree_add_69_2_groupi_n_650 & n_506);
 assign csa_tree_add_69_2_groupi_n_757 = ~(csa_tree_add_69_2_groupi_n_652 & csa_tree_add_69_2_groupi_n_288);
 assign csa_tree_add_69_2_groupi_n_756 = ~(csa_tree_add_69_2_groupi_n_650 & csa_tree_add_69_2_groupi_n_287);
 assign csa_tree_add_69_2_groupi_n_755 = ~(csa_tree_add_69_2_groupi_n_645 | csa_tree_add_69_2_groupi_n_374);
 assign csa_tree_add_69_2_groupi_n_754 = ~(csa_tree_add_69_2_groupi_n_646 & n_501);
 assign csa_tree_add_69_2_groupi_n_753 = ~(n_454 & csa_tree_add_69_2_groupi_n_375);
 assign csa_tree_add_69_2_groupi_n_752 = ~(csa_tree_add_69_2_groupi_n_646 & n_497);
 assign csa_tree_add_69_2_groupi_n_750 = ~(csa_tree_add_69_2_groupi_n_646 & csa_tree_add_69_2_groupi_n_290);
 assign csa_tree_add_69_2_groupi_n_749 = ~(csa_tree_add_69_2_groupi_n_645 | n_495);
 assign csa_tree_add_69_2_groupi_n_748 = ~(csa_tree_add_69_2_groupi_n_646 & ~csa_tree_add_69_2_groupi_n_365);
 assign csa_tree_add_69_2_groupi_n_747 = ~(n_454 & n_500);
 assign csa_tree_add_69_2_groupi_n_746 = ~(n_454 & csa_tree_add_69_2_groupi_n_381);
 assign csa_tree_add_69_2_groupi_n_745 = ~(csa_tree_add_69_2_groupi_n_646 & csa_tree_add_69_2_groupi_n_284);
 assign csa_tree_add_69_2_groupi_n_744 = ~(csa_tree_add_69_2_groupi_n_92 & csa_tree_add_69_2_groupi_n_411);
 assign csa_tree_add_69_2_groupi_n_743 = ~(csa_tree_add_69_2_groupi_n_642 & ~n_480);
 assign csa_tree_add_69_2_groupi_n_742 = ~(csa_tree_add_69_2_groupi_n_92 & n_493);
 assign csa_tree_add_69_2_groupi_n_741 = ~(csa_tree_add_69_2_groupi_n_92 & csa_tree_add_69_2_groupi_n_291);
 assign csa_tree_add_69_2_groupi_n_740 = ~(n_456 | csa_tree_add_69_2_groupi_n_397);
 assign csa_tree_add_69_2_groupi_n_739 = ~(csa_tree_add_69_2_groupi_n_644 & n_463);
 assign csa_tree_add_69_2_groupi_n_738 = ~(csa_tree_add_69_2_groupi_n_644 & n_474);
 assign csa_tree_add_69_2_groupi_n_737 = ~(csa_tree_add_69_2_groupi_n_644 & n_473);
 assign csa_tree_add_69_2_groupi_n_736 = ~(csa_tree_add_69_2_groupi_n_644 & n_475);
 assign csa_tree_add_69_2_groupi_n_772 = ~(csa_tree_add_69_2_groupi_n_585 & csa_tree_add_69_2_groupi_n_279);
 assign csa_tree_add_69_2_groupi_n_735 = ~(csa_tree_add_69_2_groupi_n_584 & csa_tree_add_69_2_groupi_n_280);
 assign csa_tree_add_69_2_groupi_n_734 = ~(({in4[0]} & csa_tree_add_69_2_groupi_n_65) | ((csa_tree_add_69_2_groupi_n_65
    & csa_tree_add_69_2_groupi_n_133) | (csa_tree_add_69_2_groupi_n_133 & {in4[0]})));
 assign csa_tree_add_69_2_groupi_n_733 = ~(csa_tree_add_69_2_groupi_n_278 | (csa_tree_add_69_2_groupi_n_256
    & csa_tree_add_69_2_groupi_n_100));
 assign csa_tree_add_69_2_groupi_n_770 = ~(csa_tree_add_69_2_groupi_n_583 & csa_tree_add_69_2_groupi_n_258);
 assign csa_tree_add_69_2_groupi_n_732 = ~(csa_tree_add_69_2_groupi_n_582 & csa_tree_add_69_2_groupi_n_276);
 assign csa_tree_add_69_2_groupi_n_731 = ~((csa_tree_add_69_2_groupi_n_573 & {in4[22]}) | (csa_tree_add_69_2_groupi_n_84
    & {in4[23]}));
 assign csa_tree_add_69_2_groupi_n_730 = ~((csa_tree_add_69_2_groupi_n_575 & {in7[22]}) | (csa_tree_add_69_2_groupi_n_87
    & {in7[23]}));
 assign csa_tree_add_69_2_groupi_n_729 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_106)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_138));
 assign csa_tree_add_69_2_groupi_n_728 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_158)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_140));
 assign csa_tree_add_69_2_groupi_n_727 = ~(csa_tree_add_69_2_groupi_n_636 & csa_tree_add_69_2_groupi_n_564);
 assign csa_tree_add_69_2_groupi_n_726 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_154)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_111));
 assign csa_tree_add_69_2_groupi_n_725 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_123)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_139));
 assign csa_tree_add_69_2_groupi_n_724 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_152)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_156));
 assign csa_tree_add_69_2_groupi_n_723 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_145)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_123));
 assign csa_tree_add_69_2_groupi_n_722 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_105)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_145));
 assign csa_tree_add_69_2_groupi_n_721 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_142)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_119));
 assign csa_tree_add_69_2_groupi_n_720 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_102)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_152));
 assign csa_tree_add_69_2_groupi_n_719 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_120)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_103));
 assign csa_tree_add_69_2_groupi_n_718 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_140)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_149));
 assign csa_tree_add_69_2_groupi_n_717 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_157)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_155));
 assign csa_tree_add_69_2_groupi_n_713 = ~csa_tree_add_69_2_groupi_n_712;
 assign csa_tree_add_69_2_groupi_n_716 = ~((csa_tree_add_69_2_groupi_n_557 & csa_tree_add_69_2_groupi_n_533)
    | (csa_tree_add_69_2_groupi_n_433 & csa_tree_add_69_2_groupi_n_136));
 assign csa_tree_add_69_2_groupi_n_708 = ~((csa_tree_add_69_2_groupi_n_557 & csa_tree_add_69_2_groupi_n_433)
    | (csa_tree_add_69_2_groupi_n_419 & csa_tree_add_69_2_groupi_n_136));
 assign csa_tree_add_69_2_groupi_n_707 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_122)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_157));
 assign csa_tree_add_69_2_groupi_n_706 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_151)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_121));
 assign csa_tree_add_69_2_groupi_n_705 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_501)
    & (csa_tree_add_69_2_groupi_n_535 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_704 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_141)
    & (csa_tree_add_69_2_groupi_n_85 | csa_tree_add_69_2_groupi_n_104));
 assign csa_tree_add_69_2_groupi_n_703 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_535)
    & (csa_tree_add_69_2_groupi_n_534 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_702 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_121)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_116));
 assign csa_tree_add_69_2_groupi_n_701 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_534)
    & (csa_tree_add_69_2_groupi_n_532 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_700 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_148)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_143));
 assign csa_tree_add_69_2_groupi_n_699 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_517)
    & (csa_tree_add_69_2_groupi_n_501 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_698 = ~(csa_tree_add_69_2_groupi_n_544 & ~(csa_tree_add_69_2_groupi_n_557
    & n_465));
 assign csa_tree_add_69_2_groupi_n_697 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_471)
    & (csa_tree_add_69_2_groupi_n_470 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_696 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_474)
    & (csa_tree_add_69_2_groupi_n_491 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_695 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_112)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_142));
 assign csa_tree_add_69_2_groupi_n_694 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_114)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_144));
 assign csa_tree_add_69_2_groupi_n_693 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_101)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_120));
 assign csa_tree_add_69_2_groupi_n_692 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_488)
    & (csa_tree_add_69_2_groupi_n_490 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_715 = ~(csa_tree_add_69_2_groupi_n_21 | (csa_tree_add_69_2_groupi_n_557
    & csa_tree_add_69_2_groupi_n_486));
 assign csa_tree_add_69_2_groupi_n_691 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_477)
    & (csa_tree_add_69_2_groupi_n_500 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_690 = ~(csa_tree_add_69_2_groupi_n_546 & ~(csa_tree_add_69_2_groupi_n_557
    & n_466));
 assign csa_tree_add_69_2_groupi_n_689 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_149)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_148));
 assign csa_tree_add_69_2_groupi_n_688 = ~(csa_tree_add_69_2_groupi_n_547 & (csa_tree_add_69_2_groupi_n_88
    | csa_tree_add_69_2_groupi_n_476));
 assign csa_tree_add_69_2_groupi_n_687 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_470)
    & (csa_tree_add_69_2_groupi_n_473 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_714 = ~(csa_tree_add_69_2_groupi_n_621 & csa_tree_add_69_2_groupi_n_545);
 assign csa_tree_add_69_2_groupi_n_686 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_483)
    & (csa_tree_add_69_2_groupi_n_477 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_685 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_500)
    & (csa_tree_add_69_2_groupi_n_518 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_684 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_518)
    & (csa_tree_add_69_2_groupi_n_517 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_683 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_491)
    & (csa_tree_add_69_2_groupi_n_471 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_712 = ~(csa_tree_add_69_2_groupi_n_634 & csa_tree_add_69_2_groupi_n_565);
 assign csa_tree_add_69_2_groupi_n_682 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_473)
    & (csa_tree_add_69_2_groupi_n_492 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_681 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_489)
    & (csa_tree_add_69_2_groupi_n_474 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_680 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_481)
    & (csa_tree_add_69_2_groupi_n_483 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_679 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_490)
    & (csa_tree_add_69_2_groupi_n_489 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_678 = ~(csa_tree_add_69_2_groupi_n_543 & ~(csa_tree_add_69_2_groupi_n_557
    & csa_tree_add_69_2_groupi_n_478));
 assign csa_tree_add_69_2_groupi_n_677 = ~((csa_tree_add_69_2_groupi_n_88 | csa_tree_add_69_2_groupi_n_492)
    & (csa_tree_add_69_2_groupi_n_481 | csa_tree_add_69_2_groupi_n_78));
 assign csa_tree_add_69_2_groupi_n_676 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_104)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_106));
 assign csa_tree_add_69_2_groupi_n_675 = ~(csa_tree_add_69_2_groupi_n_569 & ~(csa_tree_add_69_2_groupi_n_573
    & {in4[0]}));
 assign csa_tree_add_69_2_groupi_n_674 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_156)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_101));
 assign csa_tree_add_69_2_groupi_n_673 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_109)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_112));
 assign csa_tree_add_69_2_groupi_n_672 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_111)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_153));
 assign csa_tree_add_69_2_groupi_n_671 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_139)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_113));
 assign csa_tree_add_69_2_groupi_n_670 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_113)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_107));
 assign csa_tree_add_69_2_groupi_n_669 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_110)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_102));
 assign csa_tree_add_69_2_groupi_n_668 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_116)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_115));
 assign csa_tree_add_69_2_groupi_n_667 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_155)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_154));
 assign csa_tree_add_69_2_groupi_n_711 = ~(csa_tree_add_69_2_groupi_n_624 & csa_tree_add_69_2_groupi_n_542);
 assign csa_tree_add_69_2_groupi_n_666 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_115)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_122));
 assign csa_tree_add_69_2_groupi_n_665 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_107)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_114));
 assign csa_tree_add_69_2_groupi_n_710 = ~(csa_tree_add_69_2_groupi_n_620 & csa_tree_add_69_2_groupi_n_549);
 assign csa_tree_add_69_2_groupi_n_664 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_143)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_110));
 assign csa_tree_add_69_2_groupi_n_663 = ~(csa_tree_add_69_2_groupi_n_622 & csa_tree_add_69_2_groupi_n_548);
 assign csa_tree_add_69_2_groupi_n_662 = ~(csa_tree_add_69_2_groupi_n_623 & csa_tree_add_69_2_groupi_n_550);
 assign csa_tree_add_69_2_groupi_n_661 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_138)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_158));
 assign csa_tree_add_69_2_groupi_n_709 = ~(csa_tree_add_69_2_groupi_n_625 & ~(n_472 & csa_tree_add_69_2_groupi_n_136));
 assign csa_tree_add_69_2_groupi_n_660 = ~(csa_tree_add_69_2_groupi_n_638 & csa_tree_add_69_2_groupi_n_568);
 assign csa_tree_add_69_2_groupi_n_659 = ~(csa_tree_add_69_2_groupi_n_637 & csa_tree_add_69_2_groupi_n_566);
 assign csa_tree_add_69_2_groupi_n_658 = ~(csa_tree_add_69_2_groupi_n_567 & ~(csa_tree_add_69_2_groupi_n_573
    & {in4[2]}));
 assign csa_tree_add_69_2_groupi_n_657 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_144)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_151));
 assign csa_tree_add_69_2_groupi_n_656 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_118)
    & (csa_tree_add_69_2_groupi_n_82 | csa_tree_add_69_2_groupi_n_150));
 assign csa_tree_add_69_2_groupi_n_655 = ~((csa_tree_add_69_2_groupi_n_574 | csa_tree_add_69_2_groupi_n_103)
    & (csa_tree_add_69_2_groupi_n_86 | csa_tree_add_69_2_groupi_n_109));
 assign csa_tree_add_69_2_groupi_n_654 = ~((csa_tree_add_69_2_groupi_n_572 | csa_tree_add_69_2_groupi_n_150)
    & (csa_tree_add_69_2_groupi_n_83 | csa_tree_add_69_2_groupi_n_105));
 assign csa_tree_add_69_2_groupi_n_651 = ~csa_tree_add_69_2_groupi_n_652;
 assign csa_tree_add_69_2_groupi_n_649 = ~csa_tree_add_69_2_groupi_n_650;
 assign csa_tree_add_69_2_groupi_n_647 = ~n_454;
 assign csa_tree_add_69_2_groupi_n_645 = ~csa_tree_add_69_2_groupi_n_646;
 assign csa_tree_add_69_2_groupi_n_643 = ~csa_tree_add_69_2_groupi_n_644;
 assign csa_tree_add_69_2_groupi_n_92 = ~n_456;
 assign csa_tree_add_69_2_groupi_n_641 = ~csa_tree_add_69_2_groupi_n_642;
 assign csa_tree_add_69_2_groupi_n_639 = ~(n_510 & ~csa_tree_add_69_2_groupi_n_578);
 assign csa_tree_add_69_2_groupi_n_638 = ~(csa_tree_add_69_2_groupi_n_573 & {in4[1]});
 assign csa_tree_add_69_2_groupi_n_637 = ~(csa_tree_add_69_2_groupi_n_575 & {in7[1]});
 assign csa_tree_add_69_2_groupi_n_636 = ~(csa_tree_add_69_2_groupi_n_575 & {in7[2]});
 assign csa_tree_add_69_2_groupi_n_635 = ~(n_505 & ~csa_tree_add_69_2_groupi_n_576);
 assign csa_tree_add_69_2_groupi_n_634 = ~(csa_tree_add_69_2_groupi_n_575 & {in7[0]});
 assign csa_tree_add_69_2_groupi_n_633 = ~(n_473 & ~n_488);
 assign csa_tree_add_69_2_groupi_n_632 = ~(n_478 & ~n_488);
 assign csa_tree_add_69_2_groupi_n_631 = ~(csa_tree_add_69_2_groupi_n_523 & ~n_488);
 assign csa_tree_add_69_2_groupi_n_630 = ~(n_482 & ~n_488);
 assign csa_tree_add_69_2_groupi_n_629 = ~(n_474 & ~n_488);
 assign csa_tree_add_69_2_groupi_n_628 = ~(n_477 & ~n_488);
 assign csa_tree_add_69_2_groupi_n_627 = ~(n_475 & ~n_488);
 assign csa_tree_add_69_2_groupi_n_626 = ~(n_463 & ~n_488);
 assign csa_tree_add_69_2_groupi_n_625 = ~(csa_tree_add_69_2_groupi_n_557 & csa_tree_add_69_2_groupi_n_294);
 assign csa_tree_add_69_2_groupi_n_624 = ~(csa_tree_add_69_2_groupi_n_557 & n_469);
 assign csa_tree_add_69_2_groupi_n_623 = ~(csa_tree_add_69_2_groupi_n_557 & n_472);
 assign csa_tree_add_69_2_groupi_n_622 = ~(csa_tree_add_69_2_groupi_n_557 & n_471);
 assign csa_tree_add_69_2_groupi_n_621 = ~(csa_tree_add_69_2_groupi_n_557 & n_467);
 assign csa_tree_add_69_2_groupi_n_620 = ~(csa_tree_add_69_2_groupi_n_557 & n_468);
 assign csa_tree_add_69_2_groupi_n_619 = ~(n_488 | csa_tree_add_69_2_groupi_n_137);
 assign csa_tree_add_69_2_groupi_n_618 = ~(n_487 | csa_tree_add_69_2_groupi_n_100);
 assign csa_tree_add_69_2_groupi_n_617 = ~(csa_tree_add_69_2_groupi_n_90 | csa_tree_add_69_2_groupi_n_100);
 assign csa_tree_add_69_2_groupi_n_616 = ~(csa_tree_add_69_2_groupi_n_578 | csa_tree_add_69_2_groupi_n_100);
 assign csa_tree_add_69_2_groupi_n_615 = ~(csa_tree_add_69_2_groupi_n_576 | csa_tree_add_69_2_groupi_n_137);
 assign csa_tree_add_69_2_groupi_n_614 = ~(csa_tree_add_69_2_groupi_n_427 & {in7[0]});
 assign csa_tree_add_69_2_groupi_n_652 = ~(n_485 | n_459);
 assign csa_tree_add_69_2_groupi_n_650 = ~(n_486 | csa_tree_add_69_2_groupi_n_416);
 assign csa_tree_add_69_2_groupi_n_646 = ~(n_457 | ~csa_tree_add_69_2_groupi_n_413);
 assign csa_tree_add_69_2_groupi_n_644 = ~(csa_tree_add_69_2_groupi_n_579 | n_458);
 assign csa_tree_add_69_2_groupi_n_642 = ~(n_490 | csa_tree_add_69_2_groupi_n_72);
 assign csa_tree_add_69_2_groupi_n_613 = ~(csa_tree_add_69_2_groupi_n_381 & ~csa_tree_add_69_2_groupi_n_577);
 assign csa_tree_add_69_2_groupi_n_612 = ~(n_502 & ~n_487);
 assign csa_tree_add_69_2_groupi_n_611 = ~(n_504 & ~csa_tree_add_69_2_groupi_n_578);
 assign csa_tree_add_69_2_groupi_n_610 = ~(n_498 & ~n_487);
 assign csa_tree_add_69_2_groupi_n_609 = ~(n_503 | ~csa_tree_add_69_2_groupi_n_427);
 assign csa_tree_add_69_2_groupi_n_608 = ~(n_491 & ~csa_tree_add_69_2_groupi_n_90);
 assign csa_tree_add_69_2_groupi_n_607 = ~(n_487 | (csa_tree_add_69_2_groupi_n_228 & csa_tree_add_69_2_groupi_n_229));
 assign csa_tree_add_69_2_groupi_n_606 = ~(n_493 & ~csa_tree_add_69_2_groupi_n_90);
 assign csa_tree_add_69_2_groupi_n_605 = ~(n_507 & ~csa_tree_add_69_2_groupi_n_576);
 assign csa_tree_add_69_2_groupi_n_604 = ~(csa_tree_add_69_2_groupi_n_411 & ~csa_tree_add_69_2_groupi_n_90);
 assign csa_tree_add_69_2_groupi_n_603 = ~(csa_tree_add_69_2_groupi_n_322 & ~csa_tree_add_69_2_groupi_n_576);
 assign csa_tree_add_69_2_groupi_n_602 = ~(n_508 & ~csa_tree_add_69_2_groupi_n_578);
 assign csa_tree_add_69_2_groupi_n_601 = ~(n_497 & ~n_487);
 assign csa_tree_add_69_2_groupi_n_600 = ~(n_500 & ~csa_tree_add_69_2_groupi_n_577);
 assign csa_tree_add_69_2_groupi_n_599 = ~(n_496 & ~csa_tree_add_69_2_groupi_n_577);
 assign csa_tree_add_69_2_groupi_n_598 = ~(n_506 & ~csa_tree_add_69_2_groupi_n_578);
 assign csa_tree_add_69_2_groupi_n_597 = ~(n_509 | ~n_485);
 assign csa_tree_add_69_2_groupi_n_596 = ~(csa_tree_add_69_2_groupi_n_365 | ~csa_tree_add_69_2_groupi_n_580);
 assign csa_tree_add_69_2_groupi_n_595 = ~(csa_tree_add_69_2_groupi_n_353 | ~csa_tree_add_69_2_groupi_n_427);
 assign csa_tree_add_69_2_groupi_n_594 = ~(csa_tree_add_69_2_groupi_n_89 & csa_tree_add_69_2_groupi_n_407);
 assign csa_tree_add_69_2_groupi_n_593 = ~(n_494 & ~csa_tree_add_69_2_groupi_n_90);
 assign csa_tree_add_69_2_groupi_n_592 = ~(n_501 & ~n_487);
 assign csa_tree_add_69_2_groupi_n_591 = ~(n_495 | ~csa_tree_add_69_2_groupi_n_580);
 assign csa_tree_add_69_2_groupi_n_590 = ~(n_512 | ~csa_tree_add_69_2_groupi_n_89);
 assign csa_tree_add_69_2_groupi_n_589 = ~(n_499 | ~csa_tree_add_69_2_groupi_n_427);
 assign csa_tree_add_69_2_groupi_n_588 = ~(csa_tree_add_69_2_groupi_n_375 & ~csa_tree_add_69_2_groupi_n_577);
 assign csa_tree_add_69_2_groupi_n_587 = ~(n_513 & ~csa_tree_add_69_2_groupi_n_90);
 assign csa_tree_add_69_2_groupi_n_586 = ~(csa_tree_add_69_2_groupi_n_382 & ~csa_tree_add_69_2_groupi_n_577);
 assign csa_tree_add_69_2_groupi_n_585 = ~(csa_tree_add_69_2_groupi_n_255 & csa_tree_add_69_2_groupi_n_137);
 assign csa_tree_add_69_2_groupi_n_584 = ~(csa_tree_add_69_2_groupi_n_254 & csa_tree_add_69_2_groupi_n_100);
 assign csa_tree_add_69_2_groupi_n_583 = ~(csa_tree_add_69_2_groupi_n_0 & csa_tree_add_69_2_groupi_n_137);
 assign csa_tree_add_69_2_groupi_n_582 = ~(csa_tree_add_69_2_groupi_n_275 & csa_tree_add_69_2_groupi_n_137);
 assign csa_tree_add_69_2_groupi_n_581 = ~((csa_tree_add_69_2_groupi_n_432 & ~csa_tree_add_69_2_groupi_n_430)
    | (csa_tree_add_69_2_groupi_n_431 & csa_tree_add_69_2_groupi_n_430));
 assign csa_tree_add_69_2_groupi_n_580 = ~n_487;
 assign csa_tree_add_69_2_groupi_n_90 = ~csa_tree_add_69_2_groupi_n_89;
 assign csa_tree_add_69_2_groupi_n_89 = ~csa_tree_add_69_2_groupi_n_425;
 assign csa_tree_add_69_2_groupi_n_579 = ~n_488;
 assign csa_tree_add_69_2_groupi_n_578 = ~n_486;
 assign csa_tree_add_69_2_groupi_n_577 = ~csa_tree_add_69_2_groupi_n_427;
 assign csa_tree_add_69_2_groupi_n_576 = ~n_485;
 assign csa_tree_add_69_2_groupi_n_574 = ~csa_tree_add_69_2_groupi_n_575;
 assign csa_tree_add_69_2_groupi_n_572 = ~csa_tree_add_69_2_groupi_n_573;
 assign csa_tree_add_69_2_groupi_n_571 = ~(n_483 & csa_tree_add_69_2_groupi_n_72);
 assign csa_tree_add_69_2_groupi_n_570 = ~(csa_tree_add_69_2_groupi_n_441 & csa_tree_add_69_2_groupi_n_72);
 assign csa_tree_add_69_2_groupi_n_569 = ~(csa_tree_add_69_2_groupi_n_84 & {in4[1]});
 assign csa_tree_add_69_2_groupi_n_568 = ~(csa_tree_add_69_2_groupi_n_84 & {in4[2]});
 assign csa_tree_add_69_2_groupi_n_567 = ~(csa_tree_add_69_2_groupi_n_84 & {in4[3]});
 assign csa_tree_add_69_2_groupi_n_566 = ~(csa_tree_add_69_2_groupi_n_87 & {in7[2]});
 assign csa_tree_add_69_2_groupi_n_565 = ~(csa_tree_add_69_2_groupi_n_87 & {in7[1]});
 assign csa_tree_add_69_2_groupi_n_564 = ~(csa_tree_add_69_2_groupi_n_87 & {in7[3]});
 assign csa_tree_add_69_2_groupi_n_563 = ~(n_460 & csa_tree_add_69_2_groupi_n_72);
 assign csa_tree_add_69_2_groupi_n_562 = ~(n_476 & csa_tree_add_69_2_groupi_n_72);
 assign csa_tree_add_69_2_groupi_n_561 = ~(csa_tree_add_69_2_groupi_n_432 & ~csa_tree_add_69_2_groupi_n_430);
 assign csa_tree_add_69_2_groupi_n_560 = ~(n_484 | csa_tree_add_69_2_groupi_n_71);
 assign csa_tree_add_69_2_groupi_n_559 = ~(csa_tree_add_69_2_groupi_n_82 | csa_tree_add_69_2_groupi_n_100);
 assign csa_tree_add_69_2_groupi_n_558 = ~(csa_tree_add_69_2_groupi_n_85 | csa_tree_add_69_2_groupi_n_137);
 assign csa_tree_add_69_2_groupi_n_575 = ~(csa_tree_add_69_2_groupi_n_87 | csa_tree_add_69_2_groupi_n_166);
 assign csa_tree_add_69_2_groupi_n_573 = ~(csa_tree_add_69_2_groupi_n_84 | csa_tree_add_69_2_groupi_n_167);
 assign csa_tree_add_69_2_groupi_n_88 = ~csa_tree_add_69_2_groupi_n_557;
 assign csa_tree_add_69_2_groupi_n_556 = ~(n_462 & csa_tree_add_69_2_groupi_n_72);
 assign csa_tree_add_69_2_groupi_n_555 = ~(n_480 | csa_tree_add_69_2_groupi_n_71);
 assign csa_tree_add_69_2_groupi_n_554 = ~(n_479 & csa_tree_add_69_2_groupi_n_72);
 assign csa_tree_add_69_2_groupi_n_553 = ~(n_461 & csa_tree_add_69_2_groupi_n_72);
 assign csa_tree_add_69_2_groupi_n_552 = ~(csa_tree_add_69_2_groupi_n_440 & csa_tree_add_69_2_groupi_n_72);
 assign csa_tree_add_69_2_groupi_n_551 = ~(csa_tree_add_69_2_groupi_n_446 & csa_tree_add_69_2_groupi_n_72);
 assign csa_tree_add_69_2_groupi_n_550 = ~(n_471 & csa_tree_add_69_2_groupi_n_136);
 assign csa_tree_add_69_2_groupi_n_549 = ~(n_467 & csa_tree_add_69_2_groupi_n_136);
 assign csa_tree_add_69_2_groupi_n_548 = ~(csa_tree_add_69_2_groupi_n_486 & csa_tree_add_69_2_groupi_n_136);
 assign csa_tree_add_69_2_groupi_n_547 = ~(n_468 & csa_tree_add_69_2_groupi_n_136);
 assign csa_tree_add_69_2_groupi_n_546 = ~(csa_tree_add_69_2_groupi_n_478 & csa_tree_add_69_2_groupi_n_136);
 assign csa_tree_add_69_2_groupi_n_545 = ~(n_466 & csa_tree_add_69_2_groupi_n_136);
 assign csa_tree_add_69_2_groupi_n_544 = ~(n_464 & csa_tree_add_69_2_groupi_n_136);
 assign csa_tree_add_69_2_groupi_n_543 = ~(n_465 & csa_tree_add_69_2_groupi_n_136);
 assign csa_tree_add_69_2_groupi_n_542 = ~(n_470 & csa_tree_add_69_2_groupi_n_136);
 assign csa_tree_add_69_2_groupi_n_557 = ~(csa_tree_add_69_2_groupi_n_285 | csa_tree_add_69_2_groupi_n_136);
 assign csa_tree_add_69_2_groupi_n_533 = ~csa_tree_add_69_2_groupi_n_532;
 assign csa_tree_add_69_2_groupi_n_506 = ~csa_tree_add_69_2_groupi_n_505;
 assign csa_tree_add_69_2_groupi_n_504 = ~csa_tree_add_69_2_groupi_n_503;
 assign csa_tree_add_69_2_groupi_n_488 = ~n_464;
 assign csa_tree_add_69_2_groupi_n_476 = ~n_470;
 assign csa_tree_add_69_2_groupi_n_454 = ~n_478;
 assign csa_tree_add_69_2_groupi_n_450 = ~n_479;
 assign csa_tree_add_69_2_groupi_n_435 = ~n_484;
 assign csa_tree_add_69_2_groupi_n_431 = ~csa_tree_add_69_2_groupi_n_432;
 assign csa_tree_add_69_2_groupi_n_86 = ~csa_tree_add_69_2_groupi_n_87;
 assign csa_tree_add_69_2_groupi_n_87 = ~csa_tree_add_69_2_groupi_n_85;
 assign csa_tree_add_69_2_groupi_n_83 = ~csa_tree_add_69_2_groupi_n_84;
 assign csa_tree_add_69_2_groupi_n_84 = ~csa_tree_add_69_2_groupi_n_82;
 assign csa_tree_add_69_2_groupi_n_422 = ~(csa_tree_add_69_2_groupi_n_94 ^ {in7[29]});
 assign csa_tree_add_69_2_groupi_n_421 = ~(csa_tree_add_69_2_groupi_n_67 ^ {in4[27]});
 assign csa_tree_add_69_2_groupi_n_420 = ~((csa_tree_add_69_2_groupi_n_76 & ~{in7[27]}) | (csa_tree_add_69_2_groupi_n_77
    & {in7[27]}));
 assign csa_tree_add_69_2_groupi_n_419 = ~((csa_tree_add_69_2_groupi_n_130 & ~{in7[31]}) | (n_434 & {in7[31]}));
 assign csa_tree_add_69_2_groupi_n_416 = ~(csa_tree_add_69_2_groupi_n_266 | csa_tree_add_69_2_groupi_n_272);
 assign csa_tree_add_69_2_groupi_n_415 = ~((csa_tree_add_69_2_groupi_n_69 | csa_tree_add_69_2_groupi_n_127)
    & ({in4[25]} | csa_tree_add_69_2_groupi_n_96));
 assign csa_tree_add_69_2_groupi_n_414 = ~((csa_tree_add_69_2_groupi_n_70 | csa_tree_add_69_2_groupi_n_126)
    & ({in7[25]} | csa_tree_add_69_2_groupi_n_64));
 assign csa_tree_add_69_2_groupi_n_541 = ~(csa_tree_add_69_2_groupi_n_94 ^ {in7[28]});
 assign csa_tree_add_69_2_groupi_n_540 = ~(csa_tree_add_69_2_groupi_n_94 ^ {in7[26]});
 assign csa_tree_add_69_2_groupi_n_538 = ~((csa_tree_add_69_2_groupi_n_133 & ~{in4[28]}) | (csa_tree_add_69_2_groupi_n_134
    & {in4[28]}));
 assign csa_tree_add_69_2_groupi_n_537 = ~(csa_tree_add_69_2_groupi_n_133 ^ {in4[26]});
 assign csa_tree_add_69_2_groupi_n_536 = ~((csa_tree_add_69_2_groupi_n_133 & ~{in4[27]}) | (csa_tree_add_69_2_groupi_n_134
    & {in4[27]}));
 assign csa_tree_add_69_2_groupi_n_535 = ~(n_434 ^ {in7[27]});
 assign csa_tree_add_69_2_groupi_n_534 = ~(n_434 ^ {in7[28]});
 assign csa_tree_add_69_2_groupi_n_532 = ~(n_434 ^ {in7[29]});
 assign csa_tree_add_69_2_groupi_n_531 = ~(csa_tree_add_69_2_groupi_n_67 ^ {in4[26]});
 assign csa_tree_add_69_2_groupi_n_530 = ~(csa_tree_add_69_2_groupi_n_94 ^ {in7[27]});
 assign csa_tree_add_69_2_groupi_n_529 = ~((csa_tree_add_69_2_groupi_n_76 & ~{in7[26]}) | (csa_tree_add_69_2_groupi_n_77
    & {in7[26]}));
 assign csa_tree_add_69_2_groupi_n_527 = ~((csa_tree_add_69_2_groupi_n_95 & {in7[14]}) | (csa_tree_add_69_2_groupi_n_152
    & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_526 = ~(csa_tree_add_69_2_groupi_n_75 ^ {in4[28]});
 assign csa_tree_add_69_2_groupi_n_525 = ~(csa_tree_add_69_2_groupi_n_75 ^ {in4[27]});
 assign csa_tree_add_69_2_groupi_n_524 = ~((csa_tree_add_69_2_groupi_n_131 & {in4[13]}) | (csa_tree_add_69_2_groupi_n_151
    & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_523 = ~((csa_tree_add_69_2_groupi_n_104 & ~csa_tree_add_69_2_groupi_n_94)
    | ({in7[4]} & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_522 = ~((csa_tree_add_69_2_groupi_n_95 & {in7[15]}) | (csa_tree_add_69_2_groupi_n_156
    & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_519 = ~((csa_tree_add_69_2_groupi_n_95 & {in7[21]}) | (csa_tree_add_69_2_groupi_n_142
    & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_518 = ~((csa_tree_add_69_2_groupi_n_130 & {in7[24]}) | (csa_tree_add_69_2_groupi_n_160
    & n_434));
 assign csa_tree_add_69_2_groupi_n_517 = ~((csa_tree_add_69_2_groupi_n_130 & {in7[25]}) | (csa_tree_add_69_2_groupi_n_126
    & n_434));
 assign csa_tree_add_69_2_groupi_n_516 = ~((csa_tree_add_69_2_groupi_n_131 & {in4[24]}) | (csa_tree_add_69_2_groupi_n_125
    & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_515 = ~((csa_tree_add_69_2_groupi_n_131 & {in4[25]}) | (csa_tree_add_69_2_groupi_n_127
    & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_514 = ~((csa_tree_add_69_2_groupi_n_95 & {in7[24]}) | (csa_tree_add_69_2_groupi_n_160
    & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_513 = ~((csa_tree_add_69_2_groupi_n_95 & {in7[25]}) | (csa_tree_add_69_2_groupi_n_126
    & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_512 = ~((csa_tree_add_69_2_groupi_n_134 & {in4[24]}) | (csa_tree_add_69_2_groupi_n_125
    & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_511 = ~((csa_tree_add_69_2_groupi_n_134 & {in4[25]}) | (csa_tree_add_69_2_groupi_n_127
    & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_510 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[25]}) | (csa_tree_add_69_2_groupi_n_126
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_509 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[25]}) | (csa_tree_add_69_2_groupi_n_127
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_508 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[24]}) | (csa_tree_add_69_2_groupi_n_125
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_507 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[24]}) | (csa_tree_add_69_2_groupi_n_160
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_505 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[24]}) | (csa_tree_add_69_2_groupi_n_160
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_503 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[24]}) | (csa_tree_add_69_2_groupi_n_125
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_502 = ~(csa_tree_add_69_2_groupi_n_75 ^ {in4[26]});
 assign csa_tree_add_69_2_groupi_n_501 = ~(n_434 ^ {in7[26]});
 assign csa_tree_add_69_2_groupi_n_500 = ~((csa_tree_add_69_2_groupi_n_130 & {in7[23]}) | (csa_tree_add_69_2_groupi_n_124
    & n_434));
 assign csa_tree_add_69_2_groupi_n_499 = ~((csa_tree_add_69_2_groupi_n_95 & {in7[23]}) | (csa_tree_add_69_2_groupi_n_124
    & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_498 = ~((csa_tree_add_69_2_groupi_n_131 & {in4[23]}) | (csa_tree_add_69_2_groupi_n_159
    & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_497 = ~((csa_tree_add_69_2_groupi_n_134 & {in4[23]}) | (csa_tree_add_69_2_groupi_n_159
    & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_496 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[23]}) | (csa_tree_add_69_2_groupi_n_124
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_495 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[23]}) | (csa_tree_add_69_2_groupi_n_159
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_494 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[23]}) | (csa_tree_add_69_2_groupi_n_124
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_493 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[23]}) | (csa_tree_add_69_2_groupi_n_159
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_492 = ~((csa_tree_add_69_2_groupi_n_130 & {in7[19]}) | (csa_tree_add_69_2_groupi_n_109
    & n_434));
 assign csa_tree_add_69_2_groupi_n_491 = ~((csa_tree_add_69_2_groupi_n_130 & {in7[15]}) | (csa_tree_add_69_2_groupi_n_156
    & n_434));
 assign csa_tree_add_69_2_groupi_n_490 = ~((csa_tree_add_69_2_groupi_n_130 & {in7[12]}) | (csa_tree_add_69_2_groupi_n_110
    & n_434));
 assign csa_tree_add_69_2_groupi_n_489 = ~((csa_tree_add_69_2_groupi_n_130 & {in7[13]}) | (csa_tree_add_69_2_groupi_n_102
    & n_434));
 assign csa_tree_add_69_2_groupi_n_486 = ~((n_434 | csa_tree_add_69_2_groupi_n_141) & ({in7[3]} | csa_tree_add_69_2_groupi_n_130));
 assign csa_tree_add_69_2_groupi_n_483 = ~((csa_tree_add_69_2_groupi_n_130 & {in7[21]}) | (csa_tree_add_69_2_groupi_n_142
    & n_434));
 assign csa_tree_add_69_2_groupi_n_481 = ~((csa_tree_add_69_2_groupi_n_130 & {in7[20]}) | (csa_tree_add_69_2_groupi_n_112
    & n_434));
 assign csa_tree_add_69_2_groupi_n_478 = ~((csa_tree_add_69_2_groupi_n_149 & ~n_434) | ({in7[9]} & n_434));
 assign csa_tree_add_69_2_groupi_n_477 = ~((csa_tree_add_69_2_groupi_n_130 & {in7[22]}) | (csa_tree_add_69_2_groupi_n_119
    & n_434));
 assign csa_tree_add_69_2_groupi_n_474 = ~((csa_tree_add_69_2_groupi_n_130 & {in7[14]}) | (csa_tree_add_69_2_groupi_n_152
    & n_434));
 assign csa_tree_add_69_2_groupi_n_473 = ~((csa_tree_add_69_2_groupi_n_130 & {in7[18]}) | (csa_tree_add_69_2_groupi_n_103
    & n_434));
 assign csa_tree_add_69_2_groupi_n_471 = ~((csa_tree_add_69_2_groupi_n_130 & {in7[16]}) | (csa_tree_add_69_2_groupi_n_101
    & n_434));
 assign csa_tree_add_69_2_groupi_n_470 = ~((csa_tree_add_69_2_groupi_n_130 & {in7[17]}) | (csa_tree_add_69_2_groupi_n_120
    & n_434));
 assign csa_tree_add_69_2_groupi_n_468 = ~((csa_tree_add_69_2_groupi_n_131 & {in4[21]}) | (csa_tree_add_69_2_groupi_n_111
    & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_466 = ~((csa_tree_add_69_2_groupi_n_95 & {in7[16]}) | (csa_tree_add_69_2_groupi_n_101
    & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_465 = ~((csa_tree_add_69_2_groupi_n_95 & {in7[12]}) | (csa_tree_add_69_2_groupi_n_110
    & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_462 = ~((csa_tree_add_69_2_groupi_n_95 & {in7[10]}) | (csa_tree_add_69_2_groupi_n_148
    & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_461 = ~((csa_tree_add_69_2_groupi_n_95 & {in7[11]}) | (csa_tree_add_69_2_groupi_n_143
    & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_460 = ~((csa_tree_add_69_2_groupi_n_131 & {in4[16]}) | (csa_tree_add_69_2_groupi_n_115
    & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_459 = ~((csa_tree_add_69_2_groupi_n_131 & {in4[20]}) | (csa_tree_add_69_2_groupi_n_154
    & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_458 = ~((csa_tree_add_69_2_groupi_n_95 & {in7[13]}) | (csa_tree_add_69_2_groupi_n_102
    & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_455 = ~((csa_tree_add_69_2_groupi_n_95 & {in7[18]}) | (csa_tree_add_69_2_groupi_n_103
    & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_452 = ~((csa_tree_add_69_2_groupi_n_131 & {in4[14]}) | (csa_tree_add_69_2_groupi_n_121
    & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_451 = ~((csa_tree_add_69_2_groupi_n_95 & {in7[22]}) | (csa_tree_add_69_2_groupi_n_119
    & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_447 = ~((csa_tree_add_69_2_groupi_n_131 & {in4[19]}) | (csa_tree_add_69_2_groupi_n_155
    & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_446 = ~((csa_tree_add_69_2_groupi_n_113 & ~csa_tree_add_69_2_groupi_n_75)
    | ({in4[9]} & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_445 = ~((csa_tree_add_69_2_groupi_n_95 & {in7[19]}) | (csa_tree_add_69_2_groupi_n_109
    & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_443 = ~((csa_tree_add_69_2_groupi_n_95 & {in7[17]}) | (csa_tree_add_69_2_groupi_n_120
    & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_441 = ~((csa_tree_add_69_2_groupi_n_75 & ~csa_tree_add_69_2_groupi_n_107)
    | (csa_tree_add_69_2_groupi_n_131 & csa_tree_add_69_2_groupi_n_107));
 assign csa_tree_add_69_2_groupi_n_440 = ~((csa_tree_add_69_2_groupi_n_105 & ~csa_tree_add_69_2_groupi_n_75)
    | ({in4[5]} & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_439 = ~((csa_tree_add_69_2_groupi_n_131 & {in4[12]}) | (csa_tree_add_69_2_groupi_n_144
    & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_437 = ~((csa_tree_add_69_2_groupi_n_131 & {in4[22]}) | (csa_tree_add_69_2_groupi_n_153
    & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_436 = ~((csa_tree_add_69_2_groupi_n_131 & {in4[17]}) | (csa_tree_add_69_2_groupi_n_122
    & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_433 = ~((csa_tree_add_69_2_groupi_n_130 & ~{in7[30]}) | (n_434 & {in7[30]}));
 assign csa_tree_add_69_2_groupi_n_432 = ~(csa_tree_add_69_2_groupi_n_75 & ~csa_tree_add_69_2_groupi_n_283);
 assign csa_tree_add_69_2_groupi_n_430 = ~(csa_tree_add_69_2_groupi_n_226 | csa_tree_add_69_2_groupi_n_130);
 assign csa_tree_add_69_2_groupi_n_85 = ~(csa_tree_add_69_2_groupi_n_277 | csa_tree_add_69_2_groupi_n_9);
 assign csa_tree_add_69_2_groupi_n_82 = ~(csa_tree_add_69_2_groupi_n_281 | csa_tree_add_69_2_groupi_n_10);
 assign csa_tree_add_69_2_groupi_n_413 = ~((csa_tree_add_69_2_groupi_n_133 & ~csa_tree_add_69_2_groupi_n_65)
    | (csa_tree_add_69_2_groupi_n_134 & csa_tree_add_69_2_groupi_n_65));
 assign csa_tree_add_69_2_groupi_n_427 = ~(csa_tree_add_69_2_groupi_n_269 & csa_tree_add_69_2_groupi_n_268);
 assign csa_tree_add_69_2_groupi_n_425 = ~(csa_tree_add_69_2_groupi_n_262 | csa_tree_add_69_2_groupi_n_270);
 assign csa_tree_add_69_2_groupi_n_408 = ~csa_tree_add_69_2_groupi_n_407;
 assign csa_tree_add_69_2_groupi_n_390 = ~n_496;
 assign csa_tree_add_69_2_groupi_n_385 = ~n_498;
 assign csa_tree_add_69_2_groupi_n_383 = ~csa_tree_add_69_2_groupi_n_382;
 assign csa_tree_add_69_2_groupi_n_333 = ~n_507;
 assign csa_tree_add_69_2_groupi_n_326 = ~csa_tree_add_69_2_groupi_n_325;
 assign csa_tree_add_69_2_groupi_n_294 = ~((n_434 | csa_tree_add_69_2_groupi_n_137) & ({in7[0]} | csa_tree_add_69_2_groupi_n_130));
 assign csa_tree_add_69_2_groupi_n_292 = ~((csa_tree_add_69_2_groupi_n_137 & ~csa_tree_add_69_2_groupi_n_94)
    | ({in7[0]} & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_291 = ~((csa_tree_add_69_2_groupi_n_100 & ~csa_tree_add_69_2_groupi_n_133)
    | ({in4[0]} & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_290 = ~((csa_tree_add_69_2_groupi_n_100 & ~csa_tree_add_69_2_groupi_n_67)
    | ({in4[0]} & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_288 = ~((csa_tree_add_69_2_groupi_n_137 & ~csa_tree_add_69_2_groupi_n_70)
    | ({in7[0]} & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_287 = ~((csa_tree_add_69_2_groupi_n_100 & ~n_436) | ({in4[0]} & n_436));
 assign csa_tree_add_69_2_groupi_n_285 = ~(csa_tree_add_69_2_groupi_n_6 | csa_tree_add_69_2_groupi_n_172);
 assign csa_tree_add_69_2_groupi_n_412 = ~((csa_tree_add_69_2_groupi_n_134 & {in4[11]}) | (csa_tree_add_69_2_groupi_n_114
    & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_411 = ~((csa_tree_add_69_2_groupi_n_118 & ~csa_tree_add_69_2_groupi_n_133)
    | ({in4[3]} & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_410 = ~((csa_tree_add_69_2_groupi_n_134 & {in4[13]}) | (csa_tree_add_69_2_groupi_n_151
    & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_409 = ~((csa_tree_add_69_2_groupi_n_134 & {in4[15]}) | (csa_tree_add_69_2_groupi_n_116
    & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_407 = ~((csa_tree_add_69_2_groupi_n_133 | csa_tree_add_69_2_groupi_n_113)
    & ({in4[9]} | csa_tree_add_69_2_groupi_n_134));
 assign csa_tree_add_69_2_groupi_n_405 = ~((csa_tree_add_69_2_groupi_n_134 & {in4[21]}) | (csa_tree_add_69_2_groupi_n_111
    & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_404 = ~((csa_tree_add_69_2_groupi_n_134 & {in4[22]}) | (csa_tree_add_69_2_groupi_n_153
    & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_401 = ~((csa_tree_add_69_2_groupi_n_134 & {in4[19]}) | (csa_tree_add_69_2_groupi_n_155
    & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_400 = ~((csa_tree_add_69_2_groupi_n_134 & {in4[18]}) | (csa_tree_add_69_2_groupi_n_157
    & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_398 = ~((csa_tree_add_69_2_groupi_n_134 & {in4[20]}) | (csa_tree_add_69_2_groupi_n_154
    & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_397 = ~(({in4[1]} & ~n_439) | (csa_tree_add_69_2_groupi_n_108 & n_439));
 assign csa_tree_add_69_2_groupi_n_396 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[11]}) | (csa_tree_add_69_2_groupi_n_143
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_394 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[10]}) | (csa_tree_add_69_2_groupi_n_148
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_393 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[18]}) | (csa_tree_add_69_2_groupi_n_157
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_392 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[12]}) | (csa_tree_add_69_2_groupi_n_144
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_391 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[10]}) | (csa_tree_add_69_2_groupi_n_107
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_388 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[9]}) | (csa_tree_add_69_2_groupi_n_149
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_387 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[9]}) | (csa_tree_add_69_2_groupi_n_113
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_382 = ~(csa_tree_add_69_2_groupi_n_182 & ~(csa_tree_add_69_2_groupi_n_140
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_381 = ~((csa_tree_add_69_2_groupi_n_146 & ~n_382) | ({in7[1]} & n_382));
 assign csa_tree_add_69_2_groupi_n_380 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[18]}) | (csa_tree_add_69_2_groupi_n_103
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_379 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[13]}) | (csa_tree_add_69_2_groupi_n_151
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_378 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[22]}) | (csa_tree_add_69_2_groupi_n_153
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_377 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[16]}) | (csa_tree_add_69_2_groupi_n_115
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_376 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[17]}) | (csa_tree_add_69_2_groupi_n_120
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_375 = ~((csa_tree_add_69_2_groupi_n_158 & ~csa_tree_add_69_2_groupi_n_76)
    | ({in7[7]} & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_374 = ~(csa_tree_add_69_2_groupi_n_206 | ~({in4[2]} | csa_tree_add_69_2_groupi_n_66));
 assign csa_tree_add_69_2_groupi_n_284 = ~(csa_tree_add_69_2_groupi_n_228 & csa_tree_add_69_2_groupi_n_229);
 assign csa_tree_add_69_2_groupi_n_373 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[11]}) | (csa_tree_add_69_2_groupi_n_114
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_372 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[15]}) | (csa_tree_add_69_2_groupi_n_156
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_371 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[17]}) | (csa_tree_add_69_2_groupi_n_122
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_370 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[21]}) | (csa_tree_add_69_2_groupi_n_111
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_369 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[16]}) | (csa_tree_add_69_2_groupi_n_101
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_368 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[12]}) | (csa_tree_add_69_2_groupi_n_110
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_366 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[15]}) | (csa_tree_add_69_2_groupi_n_116
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_365 = ~(({in4[3]} & ~n_391) | (csa_tree_add_69_2_groupi_n_118 & n_391));
 assign csa_tree_add_69_2_groupi_n_364 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[21]}) | (csa_tree_add_69_2_groupi_n_142
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_363 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[20]}) | (csa_tree_add_69_2_groupi_n_154
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_362 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[19]}) | (csa_tree_add_69_2_groupi_n_155
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_359 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[22]}) | (csa_tree_add_69_2_groupi_n_119
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_358 = ~((csa_tree_add_69_2_groupi_n_95 & {in7[20]}) | (csa_tree_add_69_2_groupi_n_112
    & csa_tree_add_69_2_groupi_n_94));
 assign csa_tree_add_69_2_groupi_n_357 = ~((csa_tree_add_69_2_groupi_n_66 & {in4[14]}) | (csa_tree_add_69_2_groupi_n_121
    & csa_tree_add_69_2_groupi_n_67));
 assign csa_tree_add_69_2_groupi_n_356 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[19]}) | (csa_tree_add_69_2_groupi_n_109
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_355 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[20]}) | (csa_tree_add_69_2_groupi_n_112
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_354 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[13]}) | (csa_tree_add_69_2_groupi_n_102
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_353 = ~(({in7[5]} & ~csa_tree_add_69_2_groupi_n_76) | (csa_tree_add_69_2_groupi_n_106
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_350 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[16]}) | (csa_tree_add_69_2_groupi_n_115
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_349 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[12]}) | (csa_tree_add_69_2_groupi_n_110
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_348 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[7]}) | (csa_tree_add_69_2_groupi_n_123
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_347 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[8]}) | (csa_tree_add_69_2_groupi_n_140
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_346 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[17]}) | (csa_tree_add_69_2_groupi_n_122
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_345 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[17]}) | (csa_tree_add_69_2_groupi_n_120
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_344 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[15]}) | (csa_tree_add_69_2_groupi_n_116
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_343 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[16]}) | (csa_tree_add_69_2_groupi_n_101
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_341 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[10]}) | (csa_tree_add_69_2_groupi_n_148
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_340 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[22]}) | (csa_tree_add_69_2_groupi_n_153
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_339 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[11]}) | (csa_tree_add_69_2_groupi_n_114
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_337 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[20]}) | (csa_tree_add_69_2_groupi_n_112
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_335 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[13]}) | (csa_tree_add_69_2_groupi_n_151
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_334 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[8]}) | (csa_tree_add_69_2_groupi_n_139
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_331 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[14]}) | (csa_tree_add_69_2_groupi_n_121
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_330 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[6]}) | (csa_tree_add_69_2_groupi_n_138
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_329 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[22]}) | (csa_tree_add_69_2_groupi_n_119
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_328 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[7]}) | (csa_tree_add_69_2_groupi_n_158
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_325 = ~((csa_tree_add_69_2_groupi_n_105 & ~csa_tree_add_69_2_groupi_n_69)
    | ({in4[5]} & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_324 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[12]}) | (csa_tree_add_69_2_groupi_n_144
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_323 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[21]}) | (csa_tree_add_69_2_groupi_n_142
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_322 = ~((csa_tree_add_69_2_groupi_n_104 & ~csa_tree_add_69_2_groupi_n_70)
    | ({in7[4]} & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_321 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[13]}) | (csa_tree_add_69_2_groupi_n_102
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_319 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[20]}) | (csa_tree_add_69_2_groupi_n_154
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_318 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[19]}) | (csa_tree_add_69_2_groupi_n_109
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_317 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[19]}) | (csa_tree_add_69_2_groupi_n_155
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_316 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[6]}) | (csa_tree_add_69_2_groupi_n_145
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_315 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[18]}) | (csa_tree_add_69_2_groupi_n_157
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_313 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[9]}) | (csa_tree_add_69_2_groupi_n_113
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_312 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[15]}) | (csa_tree_add_69_2_groupi_n_156
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_310 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[18]}) | (csa_tree_add_69_2_groupi_n_103
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_309 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[21]}) | (csa_tree_add_69_2_groupi_n_111
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_308 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[9]}) | (csa_tree_add_69_2_groupi_n_149
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_307 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[11]}) | (csa_tree_add_69_2_groupi_n_143
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_306 = ~((csa_tree_add_69_2_groupi_n_96 & {in4[10]}) | (csa_tree_add_69_2_groupi_n_107
    & csa_tree_add_69_2_groupi_n_69));
 assign csa_tree_add_69_2_groupi_n_305 = ~((csa_tree_add_69_2_groupi_n_64 & {in7[14]}) | (csa_tree_add_69_2_groupi_n_152
    & csa_tree_add_69_2_groupi_n_70));
 assign csa_tree_add_69_2_groupi_n_304 = ~((csa_tree_add_69_2_groupi_n_77 & {in7[14]}) | (csa_tree_add_69_2_groupi_n_152
    & csa_tree_add_69_2_groupi_n_76));
 assign csa_tree_add_69_2_groupi_n_303 = ~((csa_tree_add_69_2_groupi_n_131 & {in4[15]}) | (csa_tree_add_69_2_groupi_n_116
    & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_302 = ~((csa_tree_add_69_2_groupi_n_131 & {in4[18]}) | (csa_tree_add_69_2_groupi_n_157
    & csa_tree_add_69_2_groupi_n_75));
 assign csa_tree_add_69_2_groupi_n_301 = ~((csa_tree_add_69_2_groupi_n_134 & {in4[12]}) | (csa_tree_add_69_2_groupi_n_144
    & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_300 = ~((csa_tree_add_69_2_groupi_n_134 & {in4[10]}) | (csa_tree_add_69_2_groupi_n_107
    & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_297 = ~((csa_tree_add_69_2_groupi_n_134 & {in4[16]}) | (csa_tree_add_69_2_groupi_n_115
    & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_296 = ~((csa_tree_add_69_2_groupi_n_134 & {in4[17]}) | (csa_tree_add_69_2_groupi_n_122
    & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_295 = ~((csa_tree_add_69_2_groupi_n_134 & {in4[14]}) | (csa_tree_add_69_2_groupi_n_121
    & csa_tree_add_69_2_groupi_n_133));
 assign csa_tree_add_69_2_groupi_n_281 = ~(csa_tree_add_69_2_groupi_n_68 | csa_tree_add_69_2_groupi_n_167);
 assign csa_tree_add_69_2_groupi_n_280 = (n_391 | csa_tree_add_69_2_groupi_n_74);
 assign csa_tree_add_69_2_groupi_n_279 = (n_382 | n_430);
 assign csa_tree_add_69_2_groupi_n_278 = ~(csa_tree_add_69_2_groupi_n_75 | csa_tree_add_69_2_groupi_n_163);
 assign csa_tree_add_69_2_groupi_n_277 = ~(csa_tree_add_69_2_groupi_n_70 | csa_tree_add_69_2_groupi_n_166);
 assign csa_tree_add_69_2_groupi_n_276 = ~(csa_tree_add_69_2_groupi_n_128 & ~n_434);
 assign csa_tree_add_69_2_groupi_n_275 = ~(n_434 & n_433);
 assign csa_tree_add_69_2_groupi_n_272 = ~(n_436 | csa_tree_add_69_2_groupi_n_73);
 assign csa_tree_add_69_2_groupi_n_270 = ~(n_440 | csa_tree_add_69_2_groupi_n_131);
 assign csa_tree_add_69_2_groupi_n_269 = ~(csa_tree_add_69_2_groupi_n_161 & ~n_432);
 assign csa_tree_add_69_2_groupi_n_268 = ~(csa_tree_add_69_2_groupi_n_80 & csa_tree_add_69_2_groupi_n_94);
 assign csa_tree_add_69_2_groupi_n_266 = ~(csa_tree_add_69_2_groupi_n_97 | ~csa_tree_add_69_2_groupi_n_129);
 assign csa_tree_add_69_2_groupi_n_262 = ~(csa_tree_add_69_2_groupi_n_75 | csa_tree_add_69_2_groupi_n_162);
 assign csa_tree_add_69_2_groupi_n_258 = ~(csa_tree_add_69_2_groupi_n_80 & ~n_432);
 assign csa_tree_add_69_2_groupi_n_256 = ~(csa_tree_add_69_2_groupi_n_75 & csa_tree_add_69_2_groupi_n_163);
 assign csa_tree_add_69_2_groupi_n_255 = ~(n_382 & n_430);
 assign csa_tree_add_69_2_groupi_n_254 = ~(n_391 & csa_tree_add_69_2_groupi_n_74);
 assign csa_tree_add_69_2_groupi_n_283 = ~(csa_tree_add_69_2_groupi_n_71 | csa_tree_add_69_2_groupi_n_100);
 assign csa_tree_add_69_2_groupi_n_229 = ~(csa_tree_add_69_2_groupi_n_67 & ~{in4[6]});
 assign csa_tree_add_69_2_groupi_n_228 = (csa_tree_add_69_2_groupi_n_67 | csa_tree_add_69_2_groupi_n_145);
 assign csa_tree_add_69_2_groupi_n_206 = ~(csa_tree_add_69_2_groupi_n_67 | csa_tree_add_69_2_groupi_n_147);
 assign csa_tree_add_69_2_groupi_n_182 = ~(csa_tree_add_69_2_groupi_n_77 & {in7[8]});
 assign csa_tree_add_69_2_groupi_n_172 = ~(n_434 | csa_tree_add_69_2_groupi_n_78);
 assign csa_tree_add_69_2_groupi_n_227 = ~(csa_tree_add_69_2_groupi_n_72 & csa_tree_add_69_2_groupi_n_75);
 assign csa_tree_add_69_2_groupi_n_226 = ~(csa_tree_add_69_2_groupi_n_78 | csa_tree_add_69_2_groupi_n_137);
 assign csa_tree_add_69_2_groupi_n_167 = ~n_388;
 assign csa_tree_add_69_2_groupi_n_166 = ~n_379;
 assign csa_tree_add_69_2_groupi_n_165 = ~n_430;
 assign csa_tree_add_69_2_groupi_n_163 = ~csa_tree_add_69_2_groupi_n_162;
 assign csa_tree_add_69_2_groupi_n_162 = ~n_440;
 assign csa_tree_add_69_2_groupi_n_161 = ~csa_tree_add_69_2_groupi_n_80;
 assign csa_tree_add_69_2_groupi_n_80 = ~n_431;
 assign csa_tree_add_69_2_groupi_n_160 = ~{in7[24]};
 assign csa_tree_add_69_2_groupi_n_159 = ~{in4[23]};
 assign csa_tree_add_69_2_groupi_n_158 = ~{in7[7]};
 assign csa_tree_add_69_2_groupi_n_157 = ~{in4[18]};
 assign csa_tree_add_69_2_groupi_n_156 = ~{in7[15]};
 assign csa_tree_add_69_2_groupi_n_155 = ~{in4[19]};
 assign csa_tree_add_69_2_groupi_n_154 = ~{in4[20]};
 assign csa_tree_add_69_2_groupi_n_153 = ~{in4[22]};
 assign csa_tree_add_69_2_groupi_n_152 = ~{in7[14]};
 assign csa_tree_add_69_2_groupi_n_151 = ~{in4[13]};
 assign csa_tree_add_69_2_groupi_n_150 = ~{in4[4]};
 assign csa_tree_add_69_2_groupi_n_149 = ~{in7[9]};
 assign csa_tree_add_69_2_groupi_n_148 = ~{in7[10]};
 assign csa_tree_add_69_2_groupi_n_147 = ~{in4[2]};
 assign csa_tree_add_69_2_groupi_n_146 = ~{in7[1]};
 assign csa_tree_add_69_2_groupi_n_145 = ~{in4[6]};
 assign csa_tree_add_69_2_groupi_n_144 = ~{in4[12]};
 assign csa_tree_add_69_2_groupi_n_143 = ~{in7[11]};
 assign csa_tree_add_69_2_groupi_n_142 = ~{in7[21]};
 assign csa_tree_add_69_2_groupi_n_141 = ~{in7[3]};
 assign csa_tree_add_69_2_groupi_n_140 = ~{in7[8]};
 assign csa_tree_add_69_2_groupi_n_139 = ~{in4[8]};
 assign csa_tree_add_69_2_groupi_n_138 = ~{in7[6]};
 assign csa_tree_add_69_2_groupi_n_137 = ~{in7[0]};
 assign csa_tree_add_69_2_groupi_n_136 = ~csa_tree_add_69_2_groupi_n_78;
 assign csa_tree_add_69_2_groupi_n_78 = ~n_435;
 assign csa_tree_add_69_2_groupi_n_76 = ~csa_tree_add_69_2_groupi_n_77;
 assign csa_tree_add_69_2_groupi_n_77 = ~n_382;
 assign csa_tree_add_69_2_groupi_n_133 = ~csa_tree_add_69_2_groupi_n_134;
 assign csa_tree_add_69_2_groupi_n_134 = ~n_439;
 assign csa_tree_add_69_2_groupi_n_75 = ~csa_tree_add_69_2_groupi_n_131;
 assign csa_tree_add_69_2_groupi_n_131 = ~n_441;
 assign csa_tree_add_69_2_groupi_n_130 = ~n_434;
 assign csa_tree_add_69_2_groupi_n_129 = ~n_437;
 assign csa_tree_add_69_2_groupi_n_74 = ~csa_tree_add_69_2_groupi_n_73;
 assign csa_tree_add_69_2_groupi_n_73 = ~n_437;
 assign csa_tree_add_69_2_groupi_n_128 = ~n_433;
 assign csa_tree_add_69_2_groupi_n_127 = ~{in4[25]};
 assign csa_tree_add_69_2_groupi_n_126 = ~{in7[25]};
 assign csa_tree_add_69_2_groupi_n_125 = ~{in4[24]};
 assign csa_tree_add_69_2_groupi_n_124 = ~{in7[23]};
 assign csa_tree_add_69_2_groupi_n_123 = ~{in4[7]};
 assign csa_tree_add_69_2_groupi_n_122 = ~{in4[17]};
 assign csa_tree_add_69_2_groupi_n_121 = ~{in4[14]};
 assign csa_tree_add_69_2_groupi_n_120 = ~{in7[17]};
 assign csa_tree_add_69_2_groupi_n_119 = ~{in7[22]};
 assign csa_tree_add_69_2_groupi_n_118 = ~{in4[3]};
 assign csa_tree_add_69_2_groupi_n_117 = ~{in7[2]};
 assign csa_tree_add_69_2_groupi_n_116 = ~{in4[15]};
 assign csa_tree_add_69_2_groupi_n_115 = ~{in4[16]};
 assign csa_tree_add_69_2_groupi_n_114 = ~{in4[11]};
 assign csa_tree_add_69_2_groupi_n_113 = ~{in4[9]};
 assign csa_tree_add_69_2_groupi_n_112 = ~{in7[20]};
 assign csa_tree_add_69_2_groupi_n_111 = ~{in4[21]};
 assign csa_tree_add_69_2_groupi_n_110 = ~{in7[12]};
 assign csa_tree_add_69_2_groupi_n_109 = ~{in7[19]};
 assign csa_tree_add_69_2_groupi_n_108 = ~{in4[1]};
 assign csa_tree_add_69_2_groupi_n_107 = ~{in4[10]};
 assign csa_tree_add_69_2_groupi_n_106 = ~{in7[5]};
 assign csa_tree_add_69_2_groupi_n_105 = ~{in4[5]};
 assign csa_tree_add_69_2_groupi_n_104 = ~{in7[4]};
 assign csa_tree_add_69_2_groupi_n_103 = ~{in7[18]};
 assign csa_tree_add_69_2_groupi_n_102 = ~{in7[13]};
 assign csa_tree_add_69_2_groupi_n_101 = ~{in7[16]};
 assign csa_tree_add_69_2_groupi_n_100 = ~{in4[0]};
 assign csa_tree_add_69_2_groupi_n_72 = ~csa_tree_add_69_2_groupi_n_71;
 assign csa_tree_add_69_2_groupi_n_71 = ~n_442;
 assign csa_tree_add_69_2_groupi_n_64 = ~csa_tree_add_69_2_groupi_n_70;
 assign csa_tree_add_69_2_groupi_n_70 = ~csa_tree_add_69_2_groupi_n_99;
 assign csa_tree_add_69_2_groupi_n_99 = ~n_429;
 assign csa_tree_add_69_2_groupi_n_97 = ~n_436;
 assign csa_tree_add_69_2_groupi_n_69 = ~csa_tree_add_69_2_groupi_n_96;
 assign csa_tree_add_69_2_groupi_n_68 = ~csa_tree_add_69_2_groupi_n_96;
 assign csa_tree_add_69_2_groupi_n_96 = ~n_436;
 assign csa_tree_add_69_2_groupi_n_67 = ~csa_tree_add_69_2_groupi_n_66;
 assign csa_tree_add_69_2_groupi_n_66 = ~n_391;
 assign csa_tree_add_69_2_groupi_n_94 = ~csa_tree_add_69_2_groupi_n_95;
 assign csa_tree_add_69_2_groupi_n_95 = ~n_432;
 assign csa_tree_add_69_2_groupi_n_58 = (n_444 & csa_tree_add_69_2_groupi_n_1418);
 assign csa_tree_add_69_2_groupi_n_56 = (n_445 & csa_tree_add_69_2_groupi_n_1406);
 assign csa_tree_add_69_2_groupi_n_54 = ~(csa_tree_add_69_2_groupi_n_1411 ^ csa_tree_add_69_2_groupi_n_1409);
 assign csa_tree_add_69_2_groupi_n_53 = (csa_tree_add_69_2_groupi_n_1407 & csa_tree_add_69_2_groupi_n_1309);
 assign csa_tree_add_69_2_groupi_n_52 = ~(csa_tree_add_69_2_groupi_n_1357 ^ csa_tree_add_69_2_groupi_n_1287);
 assign csa_tree_add_69_2_groupi_n_51 = (n_446 & csa_tree_add_69_2_groupi_n_1310);
 assign csa_tree_add_69_2_groupi_n_50 = (csa_tree_add_69_2_groupi_n_1311 & csa_tree_add_69_2_groupi_n_1214);
 assign csa_tree_add_69_2_groupi_n_48 = ~(csa_tree_add_69_2_groupi_n_1091 ^ csa_tree_add_69_2_groupi_n_1250);
 assign csa_tree_add_69_2_groupi_n_46 = ~(csa_tree_add_69_2_groupi_n_41 | ~csa_tree_add_69_2_groupi_n_1212);
 assign csa_tree_add_69_2_groupi_n_45 = ~(csa_tree_add_69_2_groupi_n_1023 & ~csa_tree_add_69_2_groupi_n_1142);
 assign csa_tree_add_69_2_groupi_n_44 = (csa_tree_add_69_2_groupi_n_1096 ^ csa_tree_add_69_2_groupi_n_1093);
 assign csa_tree_add_69_2_groupi_n_43 = (csa_tree_add_69_2_groupi_n_1198 & csa_tree_add_69_2_groupi_n_1011);
 assign csa_tree_add_69_2_groupi_n_42 = ~(csa_tree_add_69_2_groupi_n_1086 & ~csa_tree_add_69_2_groupi_n_1025);
 assign csa_tree_add_69_2_groupi_n_41 = ~(csa_tree_add_69_2_groupi_n_1192 | ~n_447);
 assign csa_tree_add_69_2_groupi_n_40 = ~(csa_tree_add_69_2_groupi_n_1025 & ~csa_tree_add_69_2_groupi_n_1086);
 assign csa_tree_add_69_2_groupi_n_39 = ~(csa_tree_add_69_2_groupi_n_945 ^ n_449);
 assign csa_tree_add_69_2_groupi_n_38 = (csa_tree_add_69_2_groupi_n_1012 ^ csa_tree_add_69_2_groupi_n_709);
 assign csa_tree_add_69_2_groupi_n_37 = (csa_tree_add_69_2_groupi_n_1071 & csa_tree_add_69_2_groupi_n_1074);
 assign csa_tree_add_69_2_groupi_n_36 = ~(csa_tree_add_69_2_groupi_n_862 & ~csa_tree_add_69_2_groupi_n_994);
 assign csa_tree_add_69_2_groupi_n_33 = ~(csa_tree_add_69_2_groupi_n_710 | ~csa_tree_add_69_2_groupi_n_975);
 assign csa_tree_add_69_2_groupi_n_32 = ~(csa_tree_add_69_2_groupi_n_970 | ~csa_tree_add_69_2_groupi_n_969);
 assign csa_tree_add_69_2_groupi_n_31 = ~(csa_tree_add_69_2_groupi_n_869 | ~csa_tree_add_69_2_groupi_n_968);
 assign csa_tree_add_69_2_groupi_n_29 = (csa_tree_add_69_2_groupi_n_867 & csa_tree_add_69_2_groupi_n_868);
 assign csa_tree_add_69_2_groupi_n_28 = (csa_tree_add_69_2_groupi_n_866 & csa_tree_add_69_2_groupi_n_860);
 assign csa_tree_add_69_2_groupi_n_27 = ~(csa_tree_add_69_2_groupi_n_1143 | ~csa_tree_add_69_2_groupi_n_865);
 assign csa_tree_add_69_2_groupi_n_26 = ~(csa_tree_add_69_2_groupi_n_64 | (csa_tree_add_69_2_groupi_n_33
    | ~csa_tree_add_69_2_groupi_n_772));
 assign csa_tree_add_69_2_groupi_n_24 = ~(csa_tree_add_69_2_groupi_n_967 | csa_tree_add_69_2_groupi_n_711);
 assign csa_tree_add_69_2_groupi_n_23 = ~(csa_tree_add_69_2_groupi_n_975 | ~csa_tree_add_69_2_groupi_n_710);
 assign csa_tree_add_69_2_groupi_n_22 = ~(csa_tree_add_69_2_groupi_n_643 | ~csa_tree_add_69_2_groupi_n_523);
 assign csa_tree_add_69_2_groupi_n_21 = ~(csa_tree_add_69_2_groupi_n_78 | ~n_469);
 assign csa_tree_add_69_2_groupi_n_20 = (n_481 & csa_tree_add_69_2_groupi_n_579);
 assign csa_tree_add_69_2_groupi_n_19 = (n_492 & csa_tree_add_69_2_groupi_n_89);
 assign csa_tree_add_69_2_groupi_n_18 = (csa_tree_add_69_2_groupi_n_397 | csa_tree_add_69_2_groupi_n_90);
 assign csa_tree_add_69_2_groupi_n_17 = (csa_tree_add_69_2_groupi_n_374 | n_487);
 assign csa_tree_add_69_2_groupi_n_16 = ~(n_454 & ~n_499);
 assign csa_tree_add_69_2_groupi_n_15 = ~(csa_tree_add_69_2_groupi_n_353 | ~n_454);
 assign csa_tree_add_69_2_groupi_n_14 = ~(csa_tree_add_69_2_groupi_n_645 | ~n_502);
 assign csa_tree_add_69_2_groupi_n_13 = ~(n_454 & ~n_503);
 assign csa_tree_add_69_2_groupi_n_12 = (n_511 & n_485);
 assign csa_tree_add_69_2_groupi_n_11 = ~(csa_tree_add_69_2_groupi_n_92 & ~n_512);
 assign csa_tree_add_69_2_groupi_n_10 = ~(csa_tree_add_69_2_groupi_n_96 | n_388);
 assign csa_tree_add_69_2_groupi_n_9 = ~(csa_tree_add_69_2_groupi_n_99 | n_379);
 assign csa_tree_add_69_2_groupi_n_6 = ~(csa_tree_add_69_2_groupi_n_130 | n_435);
 assign csa_tree_add_69_2_groupi_n_0 = ~(csa_tree_add_69_2_groupi_n_161 & n_432);
 assign csa_tree_add_69_2_groupi_n_93 = (csa_tree_add_69_2_groupi_n_1281 ^ (csa_tree_add_69_2_groupi_n_1092
    ^ csa_tree_add_69_2_groupi_n_1288));
 assign mul_72_11_n_230 = ~(n_397 ^ n_138);
 assign mul_72_11_n_0 = ~((n_159 & ~n_397) | (mul_72_11_n_37 & n_397));
 assign n_397 = ~(n_173 ^ n_101);
 assign mul_72_11_n_408 = ~(n_398 & ~n_175);
 assign n_173 = ((n_100 & n_176) | ((n_176 & n_98) | (n_98 & n_100)));
 assign n_398 = (n_176 ^ (n_98 ^ n_100));
 assign mul_72_11_n_225 = ~(n_174 & (mul_72_11_n_55 | mul_72_11_n_37));
 assign mul_72_11_n_282 = ~((n_399 | n_138) & (mul_72_11_n_55 | n_179));
 assign mul_72_11_n_248 = ~((n_399 | n_178) & (mul_72_11_n_55 | n_133));
 assign mul_72_11_n_274 = ~((n_399 | n_139) & (mul_72_11_n_55 | n_180));
 assign n_174 = ~n_175;
 assign n_175 = ~(n_399 | n_159);
 assign n_176 = ((n_99 & n_177) | ((n_177 & n_106) | (n_106 & n_99)));
 assign n_399 = (n_177 ^ (n_106 ^ n_99));
 assign mul_72_11_n_654 = ~(mul_72_11_n_55 | ((mul_72_11_n_1 & n_159) | (n_400 & n_401)));
 assign n_177 = ((n_107 & n_181) | ((n_181 & n_114) | (n_114 & n_107)));
 assign n_400 = (n_181 ^ (n_114 ^ n_107));
 assign mul_72_11_n_221 = ~((n_401 | n_159) & (mul_72_11_n_28 | mul_72_11_n_37));
 assign mul_72_11_n_205 = ~((n_401 | n_138) & (mul_72_11_n_28 | n_179));
 assign mul_72_11_n_189 = ~((n_401 | n_133) & (mul_72_11_n_28 | n_178));
 assign mul_72_11_n_190 = ~((n_401 | n_139) & (mul_72_11_n_28 | n_180));
 assign mul_72_11_n_176 = ~((n_401 | n_135) & (mul_72_11_n_28 | n_183));
 assign mul_72_11_n_79 = ~((n_401 | n_184) & (mul_72_11_n_28 | n_136));
 assign n_181 = ((n_115 & n_182) | ((n_182 & n_112) | (n_112 & n_115)));
 assign n_401 = (n_182 ^ (n_112 ^ n_115));
 assign mul_72_11_n_669 = ~(mul_72_11_n_28 | ((n_402 & n_403) | (mul_72_11_n_3 & n_159)));
 assign n_182 = ((n_113 & n_185) | ((n_185 & n_110) | (n_110 & n_113)));
 assign n_402 = (n_185 ^ (n_110 ^ n_113));
 assign mul_72_11_n_120 = ~((n_403 | n_135) & (mul_72_11_n_49 | n_183));
 assign mul_72_11_n_139 = ~((n_403 | n_138) & (mul_72_11_n_49 | n_179));
 assign mul_72_11_n_131 = ~((n_403 | n_133) & (mul_72_11_n_49 | n_178));
 assign mul_72_11_n_130 = ~((n_403 | n_139) & (mul_72_11_n_49 | n_180));
 assign mul_72_11_n_236 = ~((n_403 | n_159) & (mul_72_11_n_49 | mul_72_11_n_37));
 assign mul_72_11_n_119 = ~((n_403 | n_136) & (mul_72_11_n_49 | n_184));
 assign mul_72_11_n_72 = ~((n_403 | n_126) & (mul_72_11_n_49 | n_196));
 assign mul_72_11_n_108 = ~((n_403 | n_137) & (mul_72_11_n_49 | n_197));
 assign mul_72_11_n_318 = ~((n_188 | n_186) & (n_157 | n_150));
 assign mul_72_11_n_309 = ~((n_194 | n_186) & (n_169 | n_150));
 assign mul_72_11_n_314 = ~((n_192 | n_186) & (n_156 | n_150));
 assign mul_72_11_n_315 = ~((n_191 | n_186) & (mul_72_11_n_38 | n_150));
 assign mul_72_11_n_295 = ~((n_190 | n_186) & (n_125 | n_150));
 assign mul_72_11_n_311 = ~((n_146 | n_186) & (mul_72_11_n_39 | n_150));
 assign mul_72_11_n_308 = ~((n_144 | n_186) & (n_195 | n_150));
 assign mul_72_11_n_303 = ~((n_142 | n_186) & (n_193 | n_150));
 assign n_186 = ~n_150;
 assign n_185 = ((n_111 & n_187) | ((n_187 & n_108) | (n_108 & n_111)));
 assign n_403 = (n_187 ^ (n_108 ^ n_111));
 assign mul_72_11_n_279 = ~((n_142 | n_132) & (n_193 | n_189));
 assign mul_72_11_n_272 = ~((n_125 | n_132) & (n_190 | n_189));
 assign mul_72_11_n_293 = ~((n_132 | n_146) & (n_189 | mul_72_11_n_39));
 assign mul_72_11_n_285 = ~((n_144 | n_132) & (n_195 | n_189));
 assign mul_72_11_n_299 = ~((n_192 | n_132) & (n_156 | n_189));
 assign mul_72_11_n_289 = ~((n_132 | n_194) & (n_189 | n_169));
 assign mul_72_11_n_306 = ~((n_188 | n_132) & (n_157 | n_189));
 assign mul_72_11_n_300 = ~((n_191 | n_132) & (mul_72_11_n_38 | n_189));
 assign mul_72_11_n_232 = ~((mul_72_11_n_44 | n_132) & (n_120 | n_189));
 assign n_198 = ~(csa_tree_add_55_2_groupi_n_207 ^ {in3[16]});
 assign n_189 = ~n_132;
 assign mul_72_11_n_559 = ~(mul_72_11_n_49 | ((n_405 & n_159) | (mul_72_11_n_62 & n_404)));
 assign csa_tree_add_55_2_groupi_n_207 = ((csa_tree_add_55_2_groupi_n_122 & n_204) | ((n_204 & {in3[15]})
    | ({in3[15]} & csa_tree_add_55_2_groupi_n_122)));
 assign n_200 = (n_204 ^ ({in3[15]} ^ csa_tree_add_55_2_groupi_n_122));
 assign n_187 = ((n_109 & n_199) | ((n_199 & n_116) | (n_116 & n_109)));
 assign n_404 = (n_199 ^ (n_116 ^ n_109));
 assign mul_72_11_n_278 = ~((n_142 | n_131) & (n_193 | n_201));
 assign mul_72_11_n_271 = ~((n_125 | n_131) & (n_190 | n_201));
 assign mul_72_11_n_367 = ~((n_120 | n_131) & (mul_72_11_n_44 | n_201));
 assign mul_72_11_n_286 = ~((n_144 | n_131) & (n_195 | n_201));
 assign mul_72_11_n_290 = ~((n_131 | n_194) & (n_201 | n_169));
 assign mul_72_11_n_305 = ~((n_188 | n_131) & (n_157 | n_201));
 assign mul_72_11_n_294 = ~((n_131 | n_146) & (n_201 | mul_72_11_n_39));
 assign mul_72_11_n_298 = ~((n_192 | n_131) & (n_156 | n_201));
 assign mul_72_11_n_301 = ~((n_191 | n_131) & (mul_72_11_n_38 | n_201));
 assign n_201 = ~n_131;
 assign n_204 = ((csa_tree_add_55_2_groupi_n_160 & n_210) | ((n_210 & csa_tree_add_55_2_groupi_n_123)
    | (csa_tree_add_55_2_groupi_n_123 & csa_tree_add_55_2_groupi_n_160)));
 assign n_203 = (n_210 ^ (csa_tree_add_55_2_groupi_n_123 ^ csa_tree_add_55_2_groupi_n_160));
 assign mul_72_11_n_99 = ~((n_405 | n_133) & (mul_72_11_n_24 | n_178));
 assign mul_72_11_n_109 = ~((n_405 | n_138) & (mul_72_11_n_24 | n_179));
 assign mul_72_11_n_73 = ~((n_405 | n_159) & (mul_72_11_n_24 | mul_72_11_n_37));
 assign mul_72_11_n_98 = ~((n_405 | n_139) & (mul_72_11_n_24 | n_180));
 assign mul_72_11_n_90 = ~((n_405 | n_135) & (mul_72_11_n_24 | n_183));
 assign mul_72_11_n_93 = ~((n_405 | n_137) & (mul_72_11_n_24 | n_197));
 assign mul_72_11_n_92 = ~((n_405 | n_126) & (mul_72_11_n_24 | n_196));
 assign mul_72_11_n_91 = ~((n_405 | n_136) & (mul_72_11_n_24 | n_184));
 assign mul_72_11_n_71 = ~((n_405 | n_206) & (mul_72_11_n_24 | n_151));
 assign mul_72_11_n_105 = ~((n_405 | n_152) & (mul_72_11_n_24 | n_207));
 assign n_199 = ((n_117 & n_202) | ((n_202 & n_123) | (n_123 & n_117)));
 assign n_405 = (n_202 ^ (n_123 ^ n_117));
 assign mul_72_11_n_347 = ~((n_142 | n_130) & (n_193 | n_205));
 assign mul_72_11_n_146 = ~((n_125 | n_130) & (n_190 | n_205));
 assign mul_72_11_n_84 = ~((n_120 | n_130) & (mul_72_11_n_44 | n_205));
 assign mul_72_11_n_361 = ~((n_130 | n_144) & (n_205 | n_195));
 assign mul_72_11_n_277 = ~((n_146 | n_130) & (mul_72_11_n_39 | n_205));
 assign mul_72_11_n_280 = ~((n_192 | n_130) & (n_156 | n_205));
 assign mul_72_11_n_267 = ~((n_194 | n_130) & (n_169 | n_205));
 assign mul_72_11_n_287 = ~((n_188 | n_130) & (n_157 | n_205));
 assign mul_72_11_n_283 = ~((n_191 | n_130) & (mul_72_11_n_38 | n_205));
 assign mul_72_11_n_81 = ~((mul_72_11_n_45 | n_130) & (n_168 | n_205));
 assign n_205 = ~n_130;
 assign mul_72_11_n_665 = ~(mul_72_11_n_24 | ((mul_72_11_n_2 & n_159) | (n_406 & n_407)));
 assign n_210 = ((csa_tree_add_55_2_groupi_n_172 & n_214) | ((n_214 & csa_tree_add_55_2_groupi_n_161)
    | (csa_tree_add_55_2_groupi_n_161 & csa_tree_add_55_2_groupi_n_172)));
 assign n_209 = (n_214 ^ (csa_tree_add_55_2_groupi_n_161 ^ csa_tree_add_55_2_groupi_n_172));
 assign n_202 = ((n_124 & n_208) | ((n_208 & n_121) | (n_121 & n_124)));
 assign n_406 = (n_208 ^ (n_121 ^ n_124));
 assign mul_72_11_n_148 = ~((n_125 | n_129) & (n_190 | n_211));
 assign mul_72_11_n_85 = ~((n_120 | n_129) & (mul_72_11_n_44 | n_211));
 assign mul_72_11_n_201 = ~((n_168 | n_129) & (mul_72_11_n_45 | n_211));
 assign mul_72_11_n_319 = ~((n_142 | n_129) & (n_193 | n_211));
 assign mul_72_11_n_350 = ~((n_129 | n_144) & (n_211 | n_195));
 assign mul_72_11_n_268 = ~((n_129 | n_194) & (n_211 | n_169));
 assign mul_72_11_n_288 = ~((n_188 | n_129) & (n_157 | n_211));
 assign mul_72_11_n_276 = ~((n_146 | n_129) & (mul_72_11_n_39 | n_211));
 assign mul_72_11_n_281 = ~((n_192 | n_129) & (n_156 | n_211));
 assign mul_72_11_n_284 = ~((n_191 | n_129) & (mul_72_11_n_38 | n_211));
 assign n_211 = ~n_129;
 assign n_214 = ((csa_tree_add_55_2_groupi_n_174 & n_221) | ((n_221 & csa_tree_add_55_2_groupi_n_173)
    | (csa_tree_add_55_2_groupi_n_173 & csa_tree_add_55_2_groupi_n_174)));
 assign n_213 = (n_221 ^ (csa_tree_add_55_2_groupi_n_173 ^ csa_tree_add_55_2_groupi_n_174));
 assign mul_72_11_n_80 = ~((n_407 | n_159) & (mul_72_11_n_47 | mul_72_11_n_37));
 assign mul_72_11_n_86 = ~((n_407 | n_138) & (mul_72_11_n_47 | n_179));
 assign mul_72_11_n_87 = ~((n_407 | n_133) & (mul_72_11_n_47 | n_178));
 assign mul_72_11_n_88 = ~((n_407 | n_139) & (mul_72_11_n_47 | n_180));
 assign mul_72_11_n_96 = ~((n_407 | n_135) & (mul_72_11_n_47 | n_183));
 assign mul_72_11_n_97 = ~((n_407 | n_136) & (mul_72_11_n_47 | n_184));
 assign mul_72_11_n_112 = ~((n_407 | n_126) & (mul_72_11_n_47 | n_196));
 assign mul_72_11_n_111 = ~((n_407 | n_137) & (mul_72_11_n_47 | n_197));
 assign mul_72_11_n_122 = ~((n_407 | n_151) & (mul_72_11_n_47 | n_206));
 assign mul_72_11_n_123 = ~((n_407 | n_152) & (mul_72_11_n_47 | n_207));
 assign mul_72_11_n_147 = ~((n_407 | n_127) & (mul_72_11_n_47 | n_216));
 assign mul_72_11_n_76 = ~((n_407 | n_128) & (mul_72_11_n_47 | n_215));
 assign n_208 = ((n_122 & n_212) | ((n_212 & n_118) | (n_118 & n_122)));
 assign n_407 = (n_212 ^ (n_118 ^ n_122));
 assign mul_72_11_n_210 = ~((n_125 | n_128) & (n_190 | n_215));
 assign mul_72_11_n_194 = ~((n_120 | n_128) & (mul_72_11_n_44 | n_215));
 assign mul_72_11_n_166 = ~((n_168 | n_128) & (mul_72_11_n_45 | n_215));
 assign mul_72_11_n_83 = ~((n_142 | n_128) & (n_193 | n_215));
 assign mul_72_11_n_107 = ~((n_144 | n_128) & (n_195 | n_215));
 assign mul_72_11_n_203 = ~((n_194 | n_128) & (n_169 | n_215));
 assign mul_72_11_n_269 = ~((n_188 | n_128) & (n_157 | n_215));
 assign mul_72_11_n_374 = ~((n_146 | n_128) & (mul_72_11_n_39 | n_215));
 assign mul_72_11_n_378 = ~((n_192 | n_128) & (n_156 | n_215));
 assign mul_72_11_n_291 = ~((n_191 | n_128) & (mul_72_11_n_38 | n_215));
 assign n_215 = ~n_128;
 assign mul_72_11_n_558 = ~(mul_72_11_n_47 | (n_217 | (mul_72_11_n_61 & n_408)));
 assign n_221 = ((csa_tree_add_55_2_groupi_n_175 & n_223) | ((n_223 & csa_tree_add_55_2_groupi_n_184)
    | (csa_tree_add_55_2_groupi_n_184 & csa_tree_add_55_2_groupi_n_175)));
 assign n_220 = (n_223 ^ (csa_tree_add_55_2_groupi_n_184 ^ csa_tree_add_55_2_groupi_n_175));
 assign mul_72_11_n_260 = ~(n_408 ^ n_168);
 assign n_212 = ((n_119 & n_167) | ((n_167 & n_105) | (n_105 & n_119)));
 assign n_408 = (n_167 ^ (n_105 ^ n_119));
 assign mul_72_11_n_211 = ~((n_125 | n_127) & (n_190 | n_216));
 assign mul_72_11_n_193 = ~((n_120 | n_127) & (mul_72_11_n_44 | n_216));
 assign mul_72_11_n_165 = ~((n_168 | n_127) & (mul_72_11_n_45 | n_216));
 assign mul_72_11_n_219 = ~((n_127 | n_142) & (n_216 | n_193));
 assign mul_72_11_n_110 = ~((n_127 | n_144) & (n_216 | n_195));
 assign mul_72_11_n_178 = ~((n_194 | n_127) & (n_169 | n_216));
 assign mul_72_11_n_270 = ~((n_188 | n_127) & (n_157 | n_216));
 assign mul_72_11_n_375 = ~((n_146 | n_127) & (mul_72_11_n_39 | n_216));
 assign mul_72_11_n_273 = ~((n_192 | n_127) & (n_156 | n_216));
 assign mul_72_11_n_360 = ~((n_191 | n_127) & (mul_72_11_n_38 | n_216));
 assign n_216 = ~n_127;
 assign n_223 = ((csa_tree_add_55_2_groupi_n_185 & n_228) | ((n_228 & csa_tree_add_55_2_groupi_n_186)
    | (csa_tree_add_55_2_groupi_n_186 & csa_tree_add_55_2_groupi_n_185)));
 assign n_222 = (n_228 ^ (csa_tree_add_55_2_groupi_n_186 ^ csa_tree_add_55_2_groupi_n_185));
 assign mul_72_11_n_77 = ~((n_168 | n_159) & (mul_72_11_n_37 | mul_72_11_n_45));
 assign mul_72_11_n_557 = ~(n_226 | (mul_72_11_n_45 | (mul_72_11_n_60 & n_171)));
 assign mul_72_11_n_237 = ~((n_168 & ~n_171) | (mul_72_11_n_45 & n_171));
 assign mul_72_11_n_142 = ~((n_168 | n_151) & (mul_72_11_n_45 | n_206));
 assign mul_72_11_n_143 = ~((n_168 | n_152) & (mul_72_11_n_45 | n_207));
 assign mul_72_11_n_129 = ~((n_168 | n_126) & (mul_72_11_n_45 | n_196));
 assign mul_72_11_n_128 = ~((n_137 | n_168) & (n_197 | mul_72_11_n_45));
 assign mul_72_11_n_113 = ~((n_168 | n_135) & (mul_72_11_n_45 | n_183));
 assign mul_72_11_n_114 = ~((n_168 | n_136) & (mul_72_11_n_45 | n_184));
 assign mul_72_11_n_102 = ~((n_133 | n_168) & (n_178 | mul_72_11_n_45));
 assign mul_72_11_n_101 = ~((n_168 | n_139) & (mul_72_11_n_45 | n_180));
 assign mul_72_11_n_94 = ~((n_168 | n_138) & (mul_72_11_n_45 | n_179));
 assign n_217 = ~(mul_72_11_n_37 | mul_72_11_n_45);
 assign mul_72_11_n_45 = ~n_168;
 assign mul_72_11_n_161 = ~((n_120 | n_151) & (mul_72_11_n_44 | n_206));
 assign mul_72_11_n_197 = ~((n_151 | n_142) & (n_206 | n_193));
 assign mul_72_11_n_182 = ~((n_151 | n_125) & (n_206 | n_190));
 assign mul_72_11_n_209 = ~((n_144 | n_151) & (n_195 | n_206));
 assign mul_72_11_n_104 = ~((n_146 | n_151) & (mul_72_11_n_39 | n_206));
 assign mul_72_11_n_159 = ~((n_188 | n_151) & (n_157 | n_206));
 assign mul_72_11_n_215 = ~((n_194 | n_151) & (n_169 | n_206));
 assign mul_72_11_n_118 = ~((n_192 | n_151) & (n_156 | n_206));
 assign mul_72_11_n_150 = ~((n_191 | n_151) & (mul_72_11_n_38 | n_206));
 assign n_219 = ((csa_tree_add_69_2_groupi_n_1542 & n_225) | ((n_225 & n_54) | (n_54 & csa_tree_add_69_2_groupi_n_1542)));
 assign n_218 = (n_225 ^ (n_54 ^ csa_tree_add_69_2_groupi_n_1542));
 assign n_206 = ~n_151;
 assign n_228 = ((csa_tree_add_55_2_groupi_n_187 & n_234) | ((n_234 & csa_tree_add_55_2_groupi_n_180)
    | (csa_tree_add_55_2_groupi_n_180 & csa_tree_add_55_2_groupi_n_187)));
 assign n_227 = (n_234 ^ (csa_tree_add_55_2_groupi_n_180 ^ csa_tree_add_55_2_groupi_n_187));
 assign mul_72_11_n_259 = ((mul_72_11_n_44 & ~n_171) | (n_120 & n_171));
 assign mul_72_11_n_181 = ~((n_152 | n_125) & (n_207 | n_190));
 assign mul_72_11_n_160 = ~((n_120 | n_152) & (mul_72_11_n_44 | n_207));
 assign mul_72_11_n_208 = ~((n_144 | n_152) & (n_195 | n_207));
 assign mul_72_11_n_198 = ~((n_152 | n_142) & (n_207 | n_193));
 assign mul_72_11_n_216 = ~((n_194 | n_152) & (n_169 | n_207));
 assign mul_72_11_n_325 = ~((n_188 | n_152) & (n_157 | n_207));
 assign mul_72_11_n_100 = ~((n_146 | n_152) & (mul_72_11_n_39 | n_207));
 assign mul_72_11_n_132 = ~((n_192 | n_152) & (n_156 | n_207));
 assign mul_72_11_n_175 = ~((n_191 | n_152) & (mul_72_11_n_38 | n_207));
 assign n_225 = ((csa_tree_add_69_2_groupi_n_1543 & n_230) | ((n_230 & csa_tree_add_69_2_groupi_n_1540)
    | (csa_tree_add_69_2_groupi_n_1540 & csa_tree_add_69_2_groupi_n_1543)));
 assign n_224 = (n_230 ^ (csa_tree_add_69_2_groupi_n_1540 ^ csa_tree_add_69_2_groupi_n_1543));
 assign n_207 = ~n_152;
 assign n_234 = ((csa_tree_add_55_2_groupi_n_181 & n_240) | ((n_240 & csa_tree_add_55_2_groupi_n_178)
    | (csa_tree_add_55_2_groupi_n_178 & csa_tree_add_55_2_groupi_n_181)));
 assign n_233 = (n_240 ^ (csa_tree_add_55_2_groupi_n_178 ^ csa_tree_add_55_2_groupi_n_181));
 assign mul_72_11_n_141 = ~((n_120 | n_126) & (mul_72_11_n_44 | n_196));
 assign mul_72_11_n_238 = ~((n_120 & ~n_172) | (mul_72_11_n_44 & n_172));
 assign mul_72_11_n_75 = ~((n_159 | n_120) & (mul_72_11_n_37 | mul_72_11_n_44));
 assign mul_72_11_n_140 = ~((n_137 | n_120) & (n_197 | mul_72_11_n_44));
 assign mul_72_11_n_116 = ~((n_120 | n_133) & (mul_72_11_n_44 | n_178));
 assign mul_72_11_n_126 = ~((n_120 | n_135) & (mul_72_11_n_44 | n_183));
 assign mul_72_11_n_127 = ~((n_136 | n_120) & (n_184 | mul_72_11_n_44));
 assign mul_72_11_n_115 = ~((n_120 | n_139) & (mul_72_11_n_44 | n_180));
 assign mul_72_11_n_103 = ~((n_120 | n_138) & (mul_72_11_n_44 | n_179));
 assign mul_72_11_n_653 = ~(n_231 | mul_72_11_n_44);
 assign n_226 = ~(mul_72_11_n_37 | mul_72_11_n_44);
 assign mul_72_11_n_44 = ~n_120;
 assign mul_72_11_n_172 = ~((n_142 | n_126) & (n_193 | n_196));
 assign mul_72_11_n_155 = ~((n_126 | n_125) & (n_196 | n_190));
 assign mul_72_11_n_185 = ~((n_144 | n_126) & (n_195 | n_196));
 assign mul_72_11_n_196 = ~((n_194 | n_126) & (n_169 | n_196));
 assign mul_72_11_n_95 = ~((n_188 | n_126) & (n_157 | n_196));
 assign mul_72_11_n_202 = ~((n_146 | n_126) & (mul_72_11_n_39 | n_196));
 assign mul_72_11_n_213 = ~((n_192 | n_126) & (n_156 | n_196));
 assign mul_72_11_n_217 = ~((n_191 | n_126) & (mul_72_11_n_38 | n_196));
 assign n_230 = ((csa_tree_add_69_2_groupi_n_1541 & n_236) | ((n_236 & csa_tree_add_69_2_groupi_n_1564)
    | (csa_tree_add_69_2_groupi_n_1564 & csa_tree_add_69_2_groupi_n_1541)));
 assign n_229 = (n_236 ^ (csa_tree_add_69_2_groupi_n_1564 ^ csa_tree_add_69_2_groupi_n_1541));
 assign n_196 = ~n_126;
 assign n_240 = ((csa_tree_add_55_2_groupi_n_179 & n_246) | ((n_246 & csa_tree_add_55_2_groupi_n_170)
    | (csa_tree_add_55_2_groupi_n_170 & csa_tree_add_55_2_groupi_n_179)));
 assign n_239 = (n_246 ^ (csa_tree_add_55_2_groupi_n_170 ^ csa_tree_add_55_2_groupi_n_179));
 assign n_231 = ~(n_237 | (n_238 & n_232));
 assign mul_72_11_n_257 = ~((n_125 | n_172) & (n_190 | n_232));
 assign n_232 = ~n_172;
 assign mul_72_11_n_171 = ~((n_137 | n_142) & (n_197 | n_193));
 assign mul_72_11_n_156 = ~((n_125 | n_137) & (n_190 | n_197));
 assign mul_72_11_n_186 = ~((n_144 | n_137) & (n_195 | n_197));
 assign mul_72_11_n_195 = ~((n_194 | n_137) & (n_169 | n_197));
 assign mul_72_11_n_89 = ~((n_188 | n_137) & (n_157 | n_197));
 assign mul_72_11_n_204 = ~((n_146 | n_137) & (mul_72_11_n_39 | n_197));
 assign mul_72_11_n_212 = ~((n_192 | n_137) & (n_156 | n_197));
 assign mul_72_11_n_218 = ~((n_191 | n_137) & (mul_72_11_n_38 | n_197));
 assign n_236 = ((csa_tree_add_69_2_groupi_n_1565 & n_242) | ((n_242 & csa_tree_add_69_2_groupi_n_1562)
    | (csa_tree_add_69_2_groupi_n_1562 & csa_tree_add_69_2_groupi_n_1565)));
 assign n_235 = (n_242 ^ (csa_tree_add_69_2_groupi_n_1562 ^ csa_tree_add_69_2_groupi_n_1565));
 assign n_197 = ~n_137;
 assign n_246 = ((csa_tree_add_55_2_groupi_n_171 & n_254) | ((n_254 & csa_tree_add_55_2_groupi_n_156)
    | (csa_tree_add_55_2_groupi_n_156 & csa_tree_add_55_2_groupi_n_171)));
 assign n_245 = (n_254 ^ (csa_tree_add_55_2_groupi_n_156 ^ csa_tree_add_55_2_groupi_n_171));
 assign mul_72_11_n_137 = ~((n_125 | n_136) & (n_190 | n_184));
 assign mul_72_11_n_239 = ~((n_125 & ~n_143) | (n_190 & n_143));
 assign mul_72_11_n_74 = ~(n_238 & ~n_237);
 assign mul_72_11_n_136 = ~((n_125 | n_135) & (n_190 | n_183));
 assign mul_72_11_n_117 = ~((n_125 | n_138) & (n_190 | n_179));
 assign mul_72_11_n_124 = ~((n_125 | n_139) & (n_190 | n_180));
 assign mul_72_11_n_125 = ~((n_125 | n_133) & (n_190 | n_178));
 assign mul_72_11_n_222 = ~((n_125 | n_249) & (n_190 | n_163));
 assign mul_72_11_n_672 = ~(n_243 | n_190);
 assign n_237 = ~(n_159 | n_125);
 assign n_238 = ~(n_159 & n_125);
 assign n_190 = ~n_125;
 assign mul_72_11_n_158 = ~((n_144 | n_136) & (n_195 | n_184));
 assign mul_72_11_n_151 = ~((n_142 | n_136) & (n_193 | n_184));
 assign mul_72_11_n_184 = ~((n_146 | n_136) & (mul_72_11_n_39 | n_184));
 assign mul_72_11_n_192 = ~((n_192 | n_136) & (n_156 | n_184));
 assign mul_72_11_n_170 = ~((n_194 | n_136) & (n_169 | n_184));
 assign mul_72_11_n_206 = ~((n_188 | n_136) & (n_157 | n_184));
 assign mul_72_11_n_199 = ~((n_191 | n_136) & (mul_72_11_n_38 | n_184));
 assign n_242 = ((csa_tree_add_69_2_groupi_n_1563 & n_248) | ((n_248 & csa_tree_add_69_2_groupi_n_1555)
    | (csa_tree_add_69_2_groupi_n_1555 & csa_tree_add_69_2_groupi_n_1563)));
 assign n_241 = (n_248 ^ (csa_tree_add_69_2_groupi_n_1555 ^ csa_tree_add_69_2_groupi_n_1563));
 assign n_184 = ~n_136;
 assign n_254 = ((n_1 & csa_tree_add_55_2_groupi_n_157) | ((csa_tree_add_55_2_groupi_n_157 & csa_tree_add_55_2_groupi_n_138)
    | (csa_tree_add_55_2_groupi_n_138 & n_1)));
 assign n_253 = (csa_tree_add_55_2_groupi_n_157 ^ (csa_tree_add_55_2_groupi_n_138 ^ n_1));
 assign n_243 = ~(n_250 | (n_251 & n_244));
 assign mul_72_11_n_256 = ~((n_193 | n_143) & (n_142 | n_244));
 assign n_244 = ~n_143;
 assign mul_72_11_n_214 = ~((n_144 | n_135) & (n_195 | n_183));
 assign mul_72_11_n_152 = ~((n_142 | n_135) & (n_193 | n_183));
 assign mul_72_11_n_183 = ~((n_146 | n_135) & (mul_72_11_n_39 | n_183));
 assign mul_72_11_n_191 = ~((n_192 | n_135) & (n_156 | n_183));
 assign mul_72_11_n_169 = ~((n_194 | n_135) & (n_169 | n_183));
 assign mul_72_11_n_207 = ~((n_188 | n_135) & (n_157 | n_183));
 assign mul_72_11_n_200 = ~((n_191 | n_135) & (mul_72_11_n_38 | n_183));
 assign n_248 = ((csa_tree_add_69_2_groupi_n_1556 & n_256) | ((n_256 & csa_tree_add_69_2_groupi_n_1560)
    | (csa_tree_add_69_2_groupi_n_1560 & csa_tree_add_69_2_groupi_n_1556)));
 assign n_247 = (n_256 ^ (csa_tree_add_69_2_groupi_n_1560 ^ csa_tree_add_69_2_groupi_n_1556));
 assign n_183 = ~n_135;
 assign n_1 = ((n_8 & csa_tree_add_55_2_groupi_n_139) | ((csa_tree_add_55_2_groupi_n_139 & csa_tree_add_55_2_groupi_n_130)
    | (csa_tree_add_55_2_groupi_n_130 & n_8)));
 assign n_0 = (csa_tree_add_55_2_groupi_n_139 ^ (csa_tree_add_55_2_groupi_n_130 ^ n_8));
 assign mul_72_11_n_320 = ~((n_142 | n_149) & (n_193 | n_6));
 assign mul_72_11_n_240 = ~((n_142 & ~n_141) | (n_193 & n_141));
 assign mul_72_11_n_82 = ~(n_251 & ~n_250);
 assign mul_72_11_n_302 = ~((n_142 | n_163) & (n_193 | n_249));
 assign mul_72_11_n_121 = ~((n_142 | n_138) & (n_193 | n_179));
 assign mul_72_11_n_134 = ~((n_142 | n_139) & (n_193 | n_180));
 assign mul_72_11_n_135 = ~((n_142 | n_133) & (n_193 | n_178));
 assign mul_72_11_n_224 = ~((n_142 | n_5) & (n_193 | n_140));
 assign mul_72_11_n_671 = ~(n_252 | n_193);
 assign n_250 = ~(n_142 | n_159);
 assign n_251 = ~(n_142 & n_159);
 assign n_193 = ~n_142;
 assign mul_72_11_n_144 = ~((n_144 | n_133) & (n_195 | n_178));
 assign mul_72_11_n_164 = ~((n_146 | n_133) & (mul_72_11_n_39 | n_178));
 assign mul_72_11_n_174 = ~((n_192 | n_133) & (n_156 | n_178));
 assign mul_72_11_n_154 = ~((n_194 | n_133) & (n_169 | n_178));
 assign mul_72_11_n_188 = ~((n_188 | n_133) & (n_157 | n_178));
 assign mul_72_11_n_179 = ~((n_191 | n_133) & (mul_72_11_n_38 | n_178));
 assign n_256 = ((csa_tree_add_69_2_groupi_n_1561 & n_4) | ((n_4 & csa_tree_add_69_2_groupi_n_1537) |
    (csa_tree_add_69_2_groupi_n_1537 & csa_tree_add_69_2_groupi_n_1561)));
 assign n_255 = (n_4 ^ (csa_tree_add_69_2_groupi_n_1537 ^ csa_tree_add_69_2_groupi_n_1561));
 assign n_178 = ~n_133;
 assign n_252 = ~(n_257 | (n_258 & mul_72_11_n_37));
 assign mul_72_11_n_548 = ~(n_2 | (mul_72_11_n_386 & mul_72_11_n_377));
 assign n_8 = ((n_19 & csa_tree_add_55_2_groupi_n_131) | ((csa_tree_add_55_2_groupi_n_131 & csa_tree_add_55_2_groupi_n_114)
    | (csa_tree_add_55_2_groupi_n_114 & n_19)));
 assign n_7 = (csa_tree_add_55_2_groupi_n_131 ^ (csa_tree_add_55_2_groupi_n_114 ^ n_19));
 assign mul_72_11_n_255 = ~(n_258 & ~n_257);
 assign n_2 = ~(mul_72_11_n_46 | ((n_9 & n_157) | (n_10 & n_188)));
 assign n_257 = ~(n_144 | n_141);
 assign n_258 = ~(n_144 & n_141);
 assign mul_72_11_n_145 = ~((n_144 | n_139) & (n_195 | n_180));
 assign mul_72_11_n_163 = ~((n_146 | n_139) & (mul_72_11_n_39 | n_180));
 assign mul_72_11_n_173 = ~((n_192 | n_139) & (n_156 | n_180));
 assign mul_72_11_n_153 = ~((n_194 | n_139) & (n_169 | n_180));
 assign mul_72_11_n_187 = ~((n_188 | n_139) & (n_157 | n_180));
 assign mul_72_11_n_180 = ~((n_191 | n_139) & (mul_72_11_n_38 | n_180));
 assign n_9 = ~n_10;
 assign n_4 = ((csa_tree_add_69_2_groupi_n_1538 & n_21) | ((n_21 & csa_tree_add_69_2_groupi_n_1535) |
    (csa_tree_add_69_2_groupi_n_1535 & csa_tree_add_69_2_groupi_n_1538)));
 assign n_3 = (n_21 ^ (csa_tree_add_69_2_groupi_n_1535 ^ csa_tree_add_69_2_groupi_n_1538));
 assign n_10 = ~(n_24 ^ n_97);
 assign mul_72_11_n_376 = ~((n_188 & ~n_22) | (n_157 & n_22));
 assign n_180 = ~n_139;
 assign n_19 = ((n_375 & csa_tree_add_55_2_groupi_n_115) | ((csa_tree_add_55_2_groupi_n_115 & csa_tree_add_55_2_groupi_n_74)
    | (csa_tree_add_55_2_groupi_n_74 & n_375)));
 assign n_18 = (csa_tree_add_55_2_groupi_n_115 ^ (csa_tree_add_55_2_groupi_n_74 ^ n_375));
 assign mul_72_11_n_336 = ~((n_144 | n_134) & (n_195 | n_15));
 assign mul_72_11_n_241 = ~((n_144 & ~n_145) | (n_195 & n_145));
 assign mul_72_11_n_554 = ~((mul_72_11_n_167 & n_158) | (mul_72_11_n_386 & n_14));
 assign mul_72_11_n_226 = ~((n_144 | n_162) & (n_195 | n_16));
 assign mul_72_11_n_307 = ~((n_144 | n_163) & (n_195 | n_249));
 assign mul_72_11_n_322 = ~((n_144 | n_149) & (n_195 | n_6));
 assign mul_72_11_n_321 = ~((n_144 | n_140) & (n_195 | n_5));
 assign mul_72_11_n_133 = ~((n_144 | n_138) & (n_195 | n_179));
 assign mul_72_11_n_70 = ~((n_144 | n_159) & (n_195 | mul_72_11_n_37));
 assign mul_72_11_n_402 = ~(n_195 | (n_23 & n_27));
 assign n_22 = ~(n_25 ^ n_170);
 assign mul_72_11_n_304 = ~((n_188 & ~n_17) | (n_157 & n_17));
 assign mul_72_11_n_247 = ~((n_191 & ~n_17) | (mul_72_11_n_38 & n_17));
 assign n_195 = ~n_144;
 assign mul_72_11_n_149 = ~((n_146 | n_138) & (mul_72_11_n_39 | n_179));
 assign n_24 = ~(n_170 & ~n_25);
 assign mul_72_11_n_157 = ~((n_192 | n_138) & (n_156 | n_179));
 assign mul_72_11_n_138 = ~((n_194 | n_138) & (n_169 | n_179));
 assign mul_72_11_n_162 = ~((n_191 | n_138) & (mul_72_11_n_38 | n_179));
 assign mul_72_11_n_167 = ~((n_157 | n_138) & (n_188 | n_179));
 assign n_21 = ((csa_tree_add_69_2_groupi_n_1536 & n_35) | ((n_35 & csa_tree_add_69_2_groupi_n_1481)
    | (csa_tree_add_69_2_groupi_n_1481 & csa_tree_add_69_2_groupi_n_1536)));
 assign n_20 = (n_35 ^ (csa_tree_add_69_2_groupi_n_1481 ^ csa_tree_add_69_2_groupi_n_1536));
 assign mul_72_11_n_678 = ~(mul_72_11_n_38 | (n_12 & n_11));
 assign n_179 = ~n_138;
 assign mul_72_11_n_362 = ~((n_188 & ~n_28) | (n_157 & n_28));
 assign n_17 = ~(n_373 ^ n_164);
 assign mul_72_11_n_364 = ~((n_191 & ~n_28) | (mul_72_11_n_38 & n_28));
 assign mul_72_11_n_556 = ~(n_371 | (n_169 | (mul_72_11_n_59 & n_166)));
 assign mul_72_11_n_619 = ~(n_368 | (n_156 | (mul_72_11_n_63 & n_155)));
 assign n_375 = ((n_62 & csa_tree_add_55_2_groupi_n_75) | ((csa_tree_add_55_2_groupi_n_75 & csa_tree_add_55_2_groupi_n_43)
    | (csa_tree_add_55_2_groupi_n_43 & n_62)));
 assign n_374 = (csa_tree_add_55_2_groupi_n_75 ^ (csa_tree_add_55_2_groupi_n_43 ^ n_62));
 assign mul_72_11_n_292 = ((n_157 & ~n_104) | (n_188 & n_104));
 assign mul_72_11_n_373 = ~((n_188 | n_160) & (n_157 | n_370));
 assign n_12 = ~(n_13 & mul_72_11_n_37);
 assign mul_72_11_n_249 = ~(n_13 & n_11);
 assign mul_72_11_n_254 = ((n_169 & ~n_145) | (n_194 & n_145));
 assign mul_72_11_n_363 = ~((n_188 & ~n_103) | (n_157 & n_103));
 assign n_25 = ~(n_164 & ~n_373);
 assign n_14 = ~((n_157 & mul_72_11_n_37) | (n_188 & n_159));
 assign mul_72_11_n_357 = ~((n_188 | n_147) & (n_157 | n_31));
 assign mul_72_11_n_358 = ~((n_188 | n_148) & (n_157 | n_33));
 assign mul_72_11_n_345 = ~((n_188 | n_162) & (n_157 | n_16));
 assign mul_72_11_n_346 = ~((n_188 | n_134) & (n_157 | n_15));
 assign mul_72_11_n_333 = ~((n_188 | n_140) & (n_157 | n_5));
 assign mul_72_11_n_334 = ~((n_188 | n_149) & (n_157 | n_6));
 assign mul_72_11_n_317 = ~((n_188 | n_163) & (n_157 | n_249));
 assign mul_72_11_n_372 = ~((n_188 | n_161) & (n_157 | n_32));
 assign mul_72_11_n_670 = ~(mul_72_11_n_39 | (n_29 & n_369));
 assign mul_72_11_n_330 = ({out1[0]} | n_157);
 assign n_23 = (n_26 | n_145);
 assign mul_72_11_n_387 = (n_158 | n_157);
 assign n_372 = ~(csa_tree_add_69_2_groupi_n_1533 ^ n_39);
 assign n_13 = ~(n_30 & n_188);
 assign n_11 = ~(n_102 & n_157);
 assign n_188 = ~n_157;
 assign mul_72_11_n_67 = ~((n_159 | n_192) & (mul_72_11_n_37 | n_156));
 assign mul_72_11_n_244 = ~((n_192 & ~n_104) | (n_156 & n_104));
 assign mul_72_11_n_359 = ~((n_191 & ~n_104) | (mul_72_11_n_38 & n_104));
 assign mul_72_11_n_68 = ~((n_146 | n_159) & (mul_72_11_n_39 | mul_72_11_n_37));
 assign mul_72_11_n_66 = ~((n_159 | n_191) & (mul_72_11_n_38 | mul_72_11_n_37));
 assign mul_72_11_n_69 = ~(n_27 & ~n_26);
 assign n_28 = ~(n_153 ^ n_165);
 assign n_51 = ((csa_tree_add_69_2_groupi_n_1488 & csa_tree_add_69_2_groupi_n_1495) | ((csa_tree_add_69_2_groupi_n_1495
    & csa_tree_add_69_2_groupi_n_1475) | (csa_tree_add_69_2_groupi_n_1475 & csa_tree_add_69_2_groupi_n_1488)));
 assign n_50 = (csa_tree_add_69_2_groupi_n_1495 ^ (csa_tree_add_69_2_groupi_n_1475 ^ csa_tree_add_69_2_groupi_n_1488));
 assign n_43 = ((csa_tree_add_69_2_groupi_n_1527 & csa_tree_add_69_2_groupi_n_1493) | ((csa_tree_add_69_2_groupi_n_1493
    & csa_tree_add_69_2_groupi_n_1479) | (csa_tree_add_69_2_groupi_n_1479 & csa_tree_add_69_2_groupi_n_1527)));
 assign n_42 = (csa_tree_add_69_2_groupi_n_1493 ^ (csa_tree_add_69_2_groupi_n_1479 ^ csa_tree_add_69_2_groupi_n_1527));
 assign n_49 = ((csa_tree_add_69_2_groupi_n_1494 & csa_tree_add_69_2_groupi_n_1528) | ((csa_tree_add_69_2_groupi_n_1528
    & csa_tree_add_69_2_groupi_n_1436) | (csa_tree_add_69_2_groupi_n_1436 & csa_tree_add_69_2_groupi_n_1494)));
 assign n_48 = (csa_tree_add_69_2_groupi_n_1528 ^ (csa_tree_add_69_2_groupi_n_1436 ^ csa_tree_add_69_2_groupi_n_1494));
 assign n_41 = ((csa_tree_add_69_2_groupi_n_1518 & csa_tree_add_69_2_groupi_n_1489) | ((csa_tree_add_69_2_groupi_n_1489
    & csa_tree_add_69_2_groupi_n_1444) | (csa_tree_add_69_2_groupi_n_1444 & csa_tree_add_69_2_groupi_n_1518)));
 assign n_40 = (csa_tree_add_69_2_groupi_n_1489 ^ (csa_tree_add_69_2_groupi_n_1444 ^ csa_tree_add_69_2_groupi_n_1518));
 assign n_47 = ((csa_tree_add_69_2_groupi_n_1498 & csa_tree_add_69_2_groupi_n_1519) | ((csa_tree_add_69_2_groupi_n_1519
    & csa_tree_add_69_2_groupi_n_1438) | (csa_tree_add_69_2_groupi_n_1438 & csa_tree_add_69_2_groupi_n_1498)));
 assign n_46 = (csa_tree_add_69_2_groupi_n_1519 ^ (csa_tree_add_69_2_groupi_n_1438 ^ csa_tree_add_69_2_groupi_n_1498));
 assign n_57 = ((csa_tree_add_69_2_groupi_n_1492 & csa_tree_add_69_2_groupi_n_1521) | ((csa_tree_add_69_2_groupi_n_1521
    & csa_tree_add_69_2_groupi_n_1477) | (csa_tree_add_69_2_groupi_n_1477 & csa_tree_add_69_2_groupi_n_1492)));
 assign n_56 = (csa_tree_add_69_2_groupi_n_1521 ^ (csa_tree_add_69_2_groupi_n_1477 ^ csa_tree_add_69_2_groupi_n_1492));
 assign n_45 = ((csa_tree_add_69_2_groupi_n_1523 & csa_tree_add_69_2_groupi_n_1526) | ((csa_tree_add_69_2_groupi_n_1526
    & csa_tree_add_69_2_groupi_n_1458) | (csa_tree_add_69_2_groupi_n_1458 & csa_tree_add_69_2_groupi_n_1523)));
 assign n_44 = (csa_tree_add_69_2_groupi_n_1526 ^ (csa_tree_add_69_2_groupi_n_1458 ^ csa_tree_add_69_2_groupi_n_1523));
 assign n_37 = ((csa_tree_add_69_2_groupi_n_1490 & csa_tree_add_69_2_groupi_n_1524) | ((csa_tree_add_69_2_groupi_n_1524
    & csa_tree_add_69_2_groupi_n_1471) | (csa_tree_add_69_2_groupi_n_1471 & csa_tree_add_69_2_groupi_n_1490)));
 assign n_36 = (csa_tree_add_69_2_groupi_n_1524 ^ (csa_tree_add_69_2_groupi_n_1471 ^ csa_tree_add_69_2_groupi_n_1490));
 assign n_53 = ((csa_tree_add_69_2_groupi_n_1509 & csa_tree_add_69_2_groupi_n_1499) | ((csa_tree_add_69_2_groupi_n_1499
    & csa_tree_add_69_2_groupi_n_1467) | (csa_tree_add_69_2_groupi_n_1467 & csa_tree_add_69_2_groupi_n_1509)));
 assign n_52 = (csa_tree_add_69_2_groupi_n_1499 ^ (csa_tree_add_69_2_groupi_n_1467 ^ csa_tree_add_69_2_groupi_n_1509));
 assign n_55 = ((csa_tree_add_69_2_groupi_n_1486 & csa_tree_add_69_2_groupi_n_1491) | ((csa_tree_add_69_2_groupi_n_1491
    & csa_tree_add_69_2_groupi_n_1469) | (csa_tree_add_69_2_groupi_n_1469 & csa_tree_add_69_2_groupi_n_1486)));
 assign n_54 = (csa_tree_add_69_2_groupi_n_1491 ^ (csa_tree_add_69_2_groupi_n_1469 ^ csa_tree_add_69_2_groupi_n_1486));
 assign n_59 = ((csa_tree_add_69_2_groupi_n_1525 & csa_tree_add_69_2_groupi_n_1510) | ((csa_tree_add_69_2_groupi_n_1510
    & csa_tree_add_69_2_groupi_n_1448) | (csa_tree_add_69_2_groupi_n_1448 & csa_tree_add_69_2_groupi_n_1525)));
 assign n_58 = (csa_tree_add_69_2_groupi_n_1510 ^ (csa_tree_add_69_2_groupi_n_1448 ^ csa_tree_add_69_2_groupi_n_1525));
 assign n_35 = ((n_443 & csa_tree_add_69_2_groupi_n_1583) | ((csa_tree_add_69_2_groupi_n_1583 & csa_tree_add_69_2_groupi_n_1522)
    | (csa_tree_add_69_2_groupi_n_1522 & n_443)));
 assign n_34 = (csa_tree_add_69_2_groupi_n_1583 ^ (csa_tree_add_69_2_groupi_n_1522 ^ n_443));
 assign n_39 = ((csa_tree_add_69_2_groupi_n_1520 & csa_tree_add_69_2_groupi_n_1517) | ((csa_tree_add_69_2_groupi_n_1517
    & csa_tree_add_69_2_groupi_n_1454) | (csa_tree_add_69_2_groupi_n_1454 & csa_tree_add_69_2_groupi_n_1520)));
 assign n_38 = (csa_tree_add_69_2_groupi_n_1517 ^ (csa_tree_add_69_2_groupi_n_1454 ^ csa_tree_add_69_2_groupi_n_1520));
 assign mul_72_11_n_335 = ((mul_72_11_n_38 & ~n_103) | (n_191 & n_103));
 assign mul_72_11_n_251 = ~(n_377 & n_369);
 assign mul_72_11_n_351 = ~((n_146 | n_147) & (mul_72_11_n_39 | n_31));
 assign mul_72_11_n_371 = ~((n_191 | n_160) & (mul_72_11_n_38 | n_370));
 assign mul_72_11_n_370 = ~((n_191 | n_161) & (mul_72_11_n_38 | n_32));
 assign mul_72_11_n_368 = ~((n_192 | n_160) & (n_156 | n_370));
 assign mul_72_11_n_369 = ~((n_192 | n_161) & (n_156 | n_32));
 assign mul_72_11_n_242 = ~((n_194 & ~n_166) | (n_169 & n_166));
 assign mul_72_11_n_245 = ~((n_192 & ~n_155) | (n_156 & n_155));
 assign mul_72_11_n_250 = ((mul_72_11_n_38 & ~n_155) | (n_191 & n_155));
 assign mul_72_11_n_246 = ~((n_191 | n_30) & (mul_72_11_n_38 | n_102));
 assign n_378 = (csa_tree_add_69_2_groupi_n_38 ^ csa_tree_add_69_2_groupi_n_653);
 assign n_29 = (n_376 | n_159);
 assign mul_72_11_n_297 = ~((n_192 & ~n_103) | (n_156 & n_103));
 assign mul_72_11_n_243 = ~((mul_72_11_n_39 & ~n_154) | (n_146 & n_154));
 assign mul_72_11_n_253 = ((mul_72_11_n_39 & ~n_166) | (n_146 & n_166));
 assign mul_72_11_n_227 = ~((n_169 | n_148) & (n_194 | n_33));
 assign mul_72_11_n_348 = ~((n_169 | n_147) & (n_194 | n_31));
 assign mul_72_11_n_231 = ~((mul_72_11_n_39 | n_160) & (n_146 | n_370));
 assign mul_72_11_n_365 = ~((mul_72_11_n_39 | n_161) & (n_146 | n_32));
 assign n_26 = ~(n_169 | mul_72_11_n_37);
 assign n_368 = ~(mul_72_11_n_38 | mul_72_11_n_37);
 assign n_371 = ~(mul_72_11_n_39 | mul_72_11_n_37);
 assign n_27 = ~(n_169 & mul_72_11_n_37);
 assign n_373 = ~(n_165 & ~n_153);
 assign mul_72_11_n_342 = ~((n_192 | n_162) & (n_156 | n_16));
 assign mul_72_11_n_340 = ~((n_146 | n_134) & (mul_72_11_n_39 | n_15));
 assign mul_72_11_n_339 = ~((n_146 | n_162) & (mul_72_11_n_39 | n_16));
 assign mul_72_11_n_354 = ~((n_192 | n_147) & (n_156 | n_31));
 assign mul_72_11_n_353 = ~((n_192 | n_148) & (n_156 | n_33));
 assign mul_72_11_n_356 = ~((n_191 | n_147) & (mul_72_11_n_38 | n_31));
 assign mul_72_11_n_355 = ~((n_191 | n_148) & (mul_72_11_n_38 | n_33));
 assign mul_72_11_n_326 = ~((n_146 | n_140) & (mul_72_11_n_39 | n_5));
 assign mul_72_11_n_327 = ~((n_146 | n_149) & (mul_72_11_n_39 | n_6));
 assign mul_72_11_n_312 = ~((n_146 | n_163) & (mul_72_11_n_39 | n_249));
 assign mul_72_11_n_337 = ~((n_194 | n_162) & (n_169 | n_16));
 assign mul_72_11_n_338 = ~((n_194 | n_134) & (n_169 | n_15));
 assign mul_72_11_n_352 = ~((n_146 | n_148) & (mul_72_11_n_39 | n_33));
 assign mul_72_11_n_341 = ~((n_192 | n_134) & (n_156 | n_15));
 assign mul_72_11_n_343 = ~((n_191 | n_134) & (mul_72_11_n_38 | n_15));
 assign mul_72_11_n_344 = ~((n_191 | n_162) & (mul_72_11_n_38 | n_16));
 assign mul_72_11_n_324 = ~((n_194 | n_140) & (n_169 | n_5));
 assign mul_72_11_n_323 = ~((n_194 | n_149) & (n_169 | n_6));
 assign mul_72_11_n_329 = ~((n_192 | n_140) & (n_156 | n_5));
 assign mul_72_11_n_328 = ~((n_192 | n_149) & (n_156 | n_6));
 assign mul_72_11_n_331 = ~((n_191 | n_140) & (mul_72_11_n_38 | n_5));
 assign mul_72_11_n_332 = ~((n_191 | n_149) & (mul_72_11_n_38 | n_6));
 assign mul_72_11_n_310 = ~((n_194 | n_163) & (n_169 | n_249));
 assign mul_72_11_n_313 = ~((n_192 | n_163) & (n_156 | n_249));
 assign mul_72_11_n_316 = ~((n_191 | n_163) & (mul_72_11_n_38 | n_249));
 assign mul_72_11_n_46 = ~n_158;
 assign mul_72_11_n_37 = ~n_159;
 assign n_376 = ~n_377;
 assign n_377 = (n_156 | n_154);
 assign n_369 = ~(n_156 & n_154);
 assign n_32 = ~n_161;
 assign n_33 = ~n_148;
 assign n_15 = ~n_134;
 assign n_249 = ~n_163;
 assign mul_72_11_n_39 = ~n_146;
 assign n_192 = ~n_156;
 assign csa_tree_add_69_2_groupi_n_653 = (csa_tree_add_69_2_groupi_n_226 & csa_tree_add_69_2_groupi_n_283);
 assign n_60 = (csa_tree_add_69_2_groupi_n_226 ^ csa_tree_add_69_2_groupi_n_283);
 assign n_62 = (csa_tree_add_55_2_groupi_n_31 & {in3[0]});
 assign n_61 = (csa_tree_add_55_2_groupi_n_31 ^ {in3[0]});
 assign n_30 = ~n_102;
 assign n_370 = ~n_160;
 assign n_31 = ~n_147;
 assign n_16 = ~n_162;
 assign n_5 = ~n_140;
 assign n_6 = ~n_149;
 assign n_194 = ~n_169;
 assign n_191 = ~mul_72_11_n_38;
 assign n_417 = ~(csa_tree_add_55_2_groupi_n_210 ^ {in3[18]});
 assign n_424 = ~(csa_tree_add_55_2_groupi_n_222 ^ {in3[24]});
 assign n_410 = ~(csa_tree_add_55_2_groupi_n_220 ^ {in3[23]});
 assign n_419 = ~(csa_tree_add_55_2_groupi_n_226 ^ {in3[26]});
 assign n_425 = ~(csa_tree_add_55_2_groupi_n_212 ^ {in3[19]});
 assign n_423 = ~(csa_tree_add_55_2_groupi_n_218 ^ {in3[22]});
 assign n_413 = ~(csa_tree_add_55_2_groupi_n_224 ^ {in3[25]});
 assign n_426 = ~(csa_tree_add_55_2_groupi_n_216 ^ {in3[21]});
 assign n_421 = ~(csa_tree_add_69_2_groupi_n_1463 ^ csa_tree_add_69_2_groupi_n_1513);
 assign n_63 = ~((csa_tree_add_55_2_groupi_n_228 & ~{in3[27]}) | (n_416 & {in3[27]}));
 assign n_420 = ~(csa_tree_add_55_2_groupi_n_214 ^ {in3[20]});
 assign n_418 = ~(csa_tree_add_69_2_groupi_n_1548 ^ csa_tree_add_69_2_groupi_n_1482);
 assign n_411 = ~(csa_tree_add_69_2_groupi_n_1360 ^ csa_tree_add_69_2_groupi_n_1294);
 assign n_412 = ~(csa_tree_add_69_2_groupi_n_1532 ^ csa_tree_add_69_2_groupi_n_1582);
 assign n_409 = ~(csa_tree_add_69_2_groupi_n_1421 ^ csa_tree_add_69_2_groupi_n_1464);
 assign n_414 = ~(csa_tree_add_69_2_groupi_n_1217 ^ csa_tree_add_69_2_groupi_n_1094);
 assign n_422 = ~(csa_tree_add_55_2_groupi_n_208 ^ {in3[17]});
 assign n_415 = ~(n_416 & {in3[27]});
 assign n_416 = ~csa_tree_add_55_2_groupi_n_228;
 assign n_428 = ~csa_tree_add_69_2_groupi_n_1514;
 assign n_427 = ~csa_tree_add_69_2_groupi_n_1420;
 assign {out1[16]} = (mul_72_11_n_1233 ^ mul_72_11_n_1175);
 assign {out1[31]} = ~(mul_72_11_n_1314 ^ mul_72_11_n_1284);
 assign mul_72_11_n_1314 = ((mul_72_11_n_1313 & mul_72_11_n_1270) | ((mul_72_11_n_1270 & mul_72_11_n_1267)
    | (mul_72_11_n_1267 & mul_72_11_n_1313)));
 assign {out1[30]} = (mul_72_11_n_1270 ^ (mul_72_11_n_1267 ^ mul_72_11_n_1313));
 assign mul_72_11_n_1313 = ~(mul_72_11_n_1277 & (mul_72_11_n_1310 | mul_72_11_n_1281));
 assign {out1[29]} = ~(mul_72_11_n_1311 ^ mul_72_11_n_1291);
 assign mul_72_11_n_1311 = ~(mul_72_11_n_1280 & ~(mul_72_11_n_1306 & mul_72_11_n_1278));
 assign mul_72_11_n_1310 = ~(mul_72_11_n_1279 | (mul_72_11_n_1306 & mul_72_11_n_1278));
 assign {out1[28]} = ~(mul_72_11_n_1306 ^ mul_72_11_n_1290);
 assign {out1[27]} = ~(mul_72_11_n_1307 ^ mul_72_11_n_1283);
 assign mul_72_11_n_1307 = ~(mul_72_11_n_1249 & (mul_72_11_n_1302 | mul_72_11_n_1256));
 assign mul_72_11_n_1306 = ~(mul_72_11_n_1303 & (mul_72_11_n_1289 & (mul_72_11_n_1263 | mul_72_11_n_1249)));
 assign {out1[26]} = ~(mul_72_11_n_1302 ^ mul_72_11_n_1266);
 assign {out1[25]} = ~(mul_72_11_n_1301 ^ mul_72_11_n_1265);
 assign mul_72_11_n_1303 = ~(mul_72_11_n_1260 | (mul_72_11_n_1296 & (mul_72_11_n_1282 & mul_72_11_n_1261)));
 assign mul_72_11_n_1302 = ~(mul_72_11_n_1275 | (mul_72_11_n_1261 & mul_72_11_n_1296));
 assign mul_72_11_n_1301 = ~(mul_72_11_n_1244 & (mul_72_11_n_1241 | mul_72_11_n_1297));
 assign {out1[24]} = ~(mul_72_11_n_1297 ^ mul_72_11_n_1253);
 assign {out1[23]} = ~(mul_72_11_n_1298 ^ mul_72_11_n_1252);
 assign mul_72_11_n_1298 = ~(mul_72_11_n_1226 & (mul_72_11_n_1228 | mul_72_11_n_1288));
 assign mul_72_11_n_1297 = ~mul_72_11_n_1296;
 assign mul_72_11_n_1296 = ~(mul_72_11_n_1293 & (mul_72_11_n_1251 | mul_72_11_n_1262));
 assign {out1[22]} = ~(mul_72_11_n_1288 ^ mul_72_11_n_1235);
 assign {out1[21]} = ~(mul_72_11_n_1287 ^ mul_72_11_n_1229);
 assign mul_72_11_n_1293 = ~(mul_72_11_n_1243 | (mul_72_11_n_1286 | (mul_72_11_n_1250 & mul_72_11_n_1234)));
 assign {out1[19]} = ~(mul_72_11_n_1276 ^ mul_72_11_n_1205);
 assign mul_72_11_n_1291 = ~(mul_72_11_n_1277 & ~mul_72_11_n_1281);
 assign mul_72_11_n_1290 = ~(mul_72_11_n_1278 & mul_72_11_n_1280);
 assign mul_72_11_n_1289 = ~(mul_72_11_n_1275 & mul_72_11_n_1282);
 assign mul_72_11_n_1288 = ~(mul_72_11_n_1234 | (mul_72_11_n_1264 & mul_72_11_n_1227));
 assign mul_72_11_n_1287 = ~(mul_72_11_n_1211 & ~(mul_72_11_n_1264 & mul_72_11_n_1203));
 assign mul_72_11_n_1286 = ~((mul_72_11_n_1226 | mul_72_11_n_1242) & (mul_72_11_n_1262 | mul_72_11_n_1224));
 assign {out1[20]} = ~(mul_72_11_n_1264 ^ mul_72_11_n_1217);
 assign mul_72_11_n_1284 = ~(mul_72_11_n_1248 ^ mul_72_11_n_1269);
 assign mul_72_11_n_1283 = (mul_72_11_n_1263 | mul_72_11_n_1260);
 assign mul_72_11_n_1282 = ~(mul_72_11_n_1263 | mul_72_11_n_1256);
 assign mul_72_11_n_1281 = ~(mul_72_11_n_1268 | mul_72_11_n_1271);
 assign mul_72_11_n_1279 = ~mul_72_11_n_1280;
 assign mul_72_11_n_1280 = ~(mul_72_11_n_1258 & mul_72_11_n_1272);
 assign mul_72_11_n_1278 = (mul_72_11_n_1258 | mul_72_11_n_1272);
 assign mul_72_11_n_1277 = ~(mul_72_11_n_1268 & mul_72_11_n_1271);
 assign mul_72_11_n_1276 = ~(mul_72_11_n_1196 & (mul_72_11_n_1194 | mul_72_11_n_1254));
 assign mul_72_11_n_1275 = ~(mul_72_11_n_1257 & (mul_72_11_n_1255 | mul_72_11_n_1244));
 assign {out1[18]} = ~(mul_72_11_n_1254 ^ mul_72_11_n_1206);
 assign {out1[17]} = ~(mul_72_11_n_1247 ^ mul_72_11_n_1158);
 assign mul_72_11_n_1271 = ((mul_72_11_n_1221 & mul_72_11_n_1209) | ((mul_72_11_n_1209 & mul_72_11_n_1165)
    | (mul_72_11_n_1165 & mul_72_11_n_1221)));
 assign mul_72_11_n_1272 = (mul_72_11_n_1209 ^ (mul_72_11_n_1165 ^ mul_72_11_n_1221));
 assign mul_72_11_n_1269 = ((mul_72_11_n_1223 & mul_72_11_n_1207) | ((mul_72_11_n_1207 & mul_72_11_n_1182)
    | (mul_72_11_n_1182 & mul_72_11_n_1223)));
 assign mul_72_11_n_1270 = (mul_72_11_n_1207 ^ (mul_72_11_n_1182 ^ mul_72_11_n_1223));
 assign mul_72_11_n_1267 = ((mul_72_11_n_1220 & mul_72_11_n_1208) | ((mul_72_11_n_1208 & mul_72_11_n_1152)
    | (mul_72_11_n_1152 & mul_72_11_n_1220)));
 assign mul_72_11_n_1268 = (mul_72_11_n_1208 ^ (mul_72_11_n_1152 ^ mul_72_11_n_1220));
 assign mul_72_11_n_1266 = ~(mul_72_11_n_1256 | ~mul_72_11_n_1249);
 assign mul_72_11_n_1265 = ~(mul_72_11_n_1257 & ~mul_72_11_n_1255);
 assign mul_72_11_n_1264 = ~(mul_72_11_n_1251 & mul_72_11_n_1224);
 assign mul_72_11_n_1263 = ~(mul_72_11_n_1238 | mul_72_11_n_1259);
 assign mul_72_11_n_1262 = ~(mul_72_11_n_1227 & mul_72_11_n_1250);
 assign mul_72_11_n_1261 = ~(mul_72_11_n_1255 | mul_72_11_n_1241);
 assign mul_72_11_n_1260 = (mul_72_11_n_1238 & mul_72_11_n_1259);
 assign mul_72_11_n_1258 = ((mul_72_11_n_1210 & mul_72_11_n_1163) | ((mul_72_11_n_1163 & mul_72_11_n_1185)
    | (mul_72_11_n_1185 & mul_72_11_n_1210)));
 assign mul_72_11_n_1259 = (mul_72_11_n_1163 ^ (mul_72_11_n_1185 ^ mul_72_11_n_1210));
 assign mul_72_11_n_1253 = ~(mul_72_11_n_1241 | ~mul_72_11_n_1244);
 assign mul_72_11_n_1252 = (mul_72_11_n_1242 | mul_72_11_n_1243);
 assign mul_72_11_n_1257 = ~(mul_72_11_n_1230 & mul_72_11_n_1246);
 assign mul_72_11_n_1256 = ~(mul_72_11_n_1245 | mul_72_11_n_1239);
 assign mul_72_11_n_1255 = ~(mul_72_11_n_1230 | mul_72_11_n_1246);
 assign mul_72_11_n_1254 = ~(mul_72_11_n_1193 | mul_72_11_n_1240);
 assign mul_72_11_n_1251 = ~(mul_72_11_n_1204 & mul_72_11_n_1240);
 assign mul_72_11_n_1248 = ~(mul_72_11_n_1232 ^ mul_72_11_n_1189);
 assign mul_72_11_n_1247 = ~(mul_72_11_n_1172 & (mul_72_11_n_1171 | mul_72_11_n_1233));
 assign mul_72_11_n_1250 = ~(mul_72_11_n_1228 | mul_72_11_n_1242);
 assign mul_72_11_n_1249 = ~(mul_72_11_n_1245 & mul_72_11_n_1239);
 assign mul_72_11_n_1245 = ((mul_72_11_n_1180 & mul_72_11_n_1177) | ((mul_72_11_n_1177 & mul_72_11_n_1156)
    | (mul_72_11_n_1156 & mul_72_11_n_1180)));
 assign mul_72_11_n_1246 = (mul_72_11_n_1177 ^ (mul_72_11_n_1156 ^ mul_72_11_n_1180));
 assign mul_72_11_n_1244 = ~(mul_72_11_n_1231 & mul_72_11_n_1236);
 assign mul_72_11_n_1243 = (mul_72_11_n_1218 & mul_72_11_n_1237);
 assign mul_72_11_n_1242 = ~(mul_72_11_n_1218 | mul_72_11_n_1237);
 assign mul_72_11_n_1241 = ~(mul_72_11_n_1231 | mul_72_11_n_1236);
 assign mul_72_11_n_1240 = ~(mul_72_11_n_1171 | (mul_72_11_n_1149 | mul_72_11_n_1233));
 assign mul_72_11_n_1238 = ((mul_72_11_n_1179 & mul_72_11_n_1186) | ((mul_72_11_n_1186 & mul_72_11_n_1155)
    | (mul_72_11_n_1155 & mul_72_11_n_1179)));
 assign mul_72_11_n_1239 = (mul_72_11_n_1186 ^ (mul_72_11_n_1155 ^ mul_72_11_n_1179));
 assign mul_72_11_n_1236 = ((mul_72_11_n_1167 & mul_72_11_n_1110) | ((mul_72_11_n_1110 & mul_72_11_n_1168)
    | (mul_72_11_n_1168 & mul_72_11_n_1167)));
 assign mul_72_11_n_1237 = (mul_72_11_n_1110 ^ (mul_72_11_n_1168 ^ mul_72_11_n_1167));
 assign mul_72_11_n_1235 = ~(mul_72_11_n_1228 | ~mul_72_11_n_1226);
 assign mul_72_11_n_1234 = ~(mul_72_11_n_1216 & (mul_72_11_n_1215 | mul_72_11_n_1211));
 assign mul_72_11_n_1233 = ~(mul_72_11_n_1225 | ~(mul_72_11_n_1197 | mul_72_11_n_1114));
 assign mul_72_11_n_1232 = ~(mul_72_11_n_1222 ^ mul_72_11_n_1181);
 assign mul_72_11_n_1230 = ((mul_72_11_n_1166 & mul_72_11_n_1178) | ((mul_72_11_n_1178 & mul_72_11_n_1127)
    | (mul_72_11_n_1127 & mul_72_11_n_1166)));
 assign mul_72_11_n_1231 = (mul_72_11_n_1178 ^ (mul_72_11_n_1127 ^ mul_72_11_n_1166));
 assign mul_72_11_n_1229 = ~(mul_72_11_n_1216 & ~mul_72_11_n_1215);
 assign mul_72_11_n_1228 = ~(mul_72_11_n_1219 | mul_72_11_n_1212);
 assign mul_72_11_n_1227 = ~(mul_72_11_n_1215 | ~mul_72_11_n_1203);
 assign mul_72_11_n_1226 = ~(mul_72_11_n_1219 & mul_72_11_n_1212);
 assign mul_72_11_n_1225 = ~(mul_72_11_n_1173 & (mul_72_11_n_1201 & (mul_72_11_n_1119 | mul_72_11_n_1197)));
 assign mul_72_11_n_1224 = ~(mul_72_11_n_1202 | (mul_72_11_n_1198 | (mul_72_11_n_1193 & mul_72_11_n_1204)));
 assign mul_72_11_n_1222 = ((mul_72_11_n_1151 & mul_72_11_n_1095) | ((mul_72_11_n_1095 & mul_72_11_n_1141)
    | (mul_72_11_n_1141 & mul_72_11_n_1151)));
 assign mul_72_11_n_1223 = (mul_72_11_n_1095 ^ (mul_72_11_n_1141 ^ mul_72_11_n_1151));
 assign mul_72_11_n_1220 = ((mul_72_11_n_1129 & mul_72_11_n_1162) | ((mul_72_11_n_1162 & mul_72_11_n_1061)
    | (mul_72_11_n_1061 & mul_72_11_n_1129)));
 assign mul_72_11_n_1221 = (mul_72_11_n_1162 ^ (mul_72_11_n_1061 ^ mul_72_11_n_1129));
 assign mul_72_11_n_1218 = ((mul_72_11_n_1122 & mul_72_11_n_1169) | ((mul_72_11_n_1169 & mul_72_11_n_1093)
    | (mul_72_11_n_1093 & mul_72_11_n_1122)));
 assign mul_72_11_n_1219 = (mul_72_11_n_1169 ^ (mul_72_11_n_1093 ^ mul_72_11_n_1122));
 assign mul_72_11_n_1217 = ~(mul_72_11_n_1203 & mul_72_11_n_1211);
 assign mul_72_11_n_1216 = ~(mul_72_11_n_1199 & mul_72_11_n_1213);
 assign mul_72_11_n_1215 = ~(mul_72_11_n_1199 | mul_72_11_n_1213);
 assign {out1[15]} = ~(mul_72_11_n_1190 ^ mul_72_11_n_1176);
 assign mul_72_11_n_1209 = ((mul_72_11_n_1142 & mul_72_11_n_1100) | ((mul_72_11_n_1100 & mul_72_11_n_1125)
    | (mul_72_11_n_1125 & mul_72_11_n_1142)));
 assign mul_72_11_n_1210 = (mul_72_11_n_1100 ^ (mul_72_11_n_1125 ^ mul_72_11_n_1142));
 assign mul_72_11_n_1212 = ((mul_72_11_n_1123 & mul_72_11_n_1084) | ((mul_72_11_n_1084 & mul_72_11_n_1130)
    | (mul_72_11_n_1130 & mul_72_11_n_1123)));
 assign mul_72_11_n_1213 = (mul_72_11_n_1084 ^ (mul_72_11_n_1130 ^ mul_72_11_n_1123));
 assign mul_72_11_n_1207 = ((mul_72_11_n_1164 & mul_72_11_n_1128) | ((mul_72_11_n_1128 & mul_72_11_n_1108)
    | (mul_72_11_n_1108 & mul_72_11_n_1164)));
 assign mul_72_11_n_1208 = (mul_72_11_n_1128 ^ (mul_72_11_n_1108 ^ mul_72_11_n_1164));
 assign mul_72_11_n_1206 = ~(mul_72_11_n_1194 | ~mul_72_11_n_1196);
 assign mul_72_11_n_1205 = (mul_72_11_n_1195 | mul_72_11_n_1198);
 assign mul_72_11_n_1211 = ~(mul_72_11_n_1187 & mul_72_11_n_1200);
 assign mul_72_11_n_1202 = ~(mul_72_11_n_1196 | mul_72_11_n_1195);
 assign mul_72_11_n_1201 = ~((mul_72_11_n_1138 & mul_72_11_n_1174) | (mul_72_11_n_1170 & mul_72_11_n_1133));
 assign mul_72_11_n_1204 = ~(mul_72_11_n_1194 | mul_72_11_n_1195);
 assign mul_72_11_n_1203 = (mul_72_11_n_1187 | mul_72_11_n_1200);
 assign mul_72_11_n_1199 = ((mul_72_11_n_1131 & mul_72_11_n_1111) | ((mul_72_11_n_1111 & mul_72_11_n_1047)
    | (mul_72_11_n_1047 & mul_72_11_n_1131)));
 assign mul_72_11_n_1200 = (mul_72_11_n_1111 ^ (mul_72_11_n_1047 ^ mul_72_11_n_1131));
 assign mul_72_11_n_1198 = (mul_72_11_n_1188 & mul_72_11_n_1183);
 assign mul_72_11_n_1197 = ~(mul_72_11_n_1120 & mul_72_11_n_1174);
 assign mul_72_11_n_1196 = ~(mul_72_11_n_1146 & mul_72_11_n_1184);
 assign mul_72_11_n_1195 = ~(mul_72_11_n_1188 | mul_72_11_n_1183);
 assign mul_72_11_n_1194 = ~(mul_72_11_n_1146 | mul_72_11_n_1184);
 assign {out1[14]} = ~(mul_72_11_n_1161 ^ mul_72_11_n_1139);
 assign {out1[13]} = ~(mul_72_11_n_1157 ^ mul_72_11_n_1121);
 assign mul_72_11_n_1190 = ~(mul_72_11_n_1132 & (mul_72_11_n_1161 | mul_72_11_n_1134));
 assign mul_72_11_n_1189 = ~(mul_72_11_n_1159 ^ mul_72_11_n_1148);
 assign mul_72_11_n_1193 = ~(mul_72_11_n_1150 & (mul_72_11_n_1172 | mul_72_11_n_1149));
 assign mul_72_11_n_1187 = ((mul_72_11_n_1112 & mul_72_11_n_1098) | ((mul_72_11_n_1098 & mul_72_11_n_1067)
    | (mul_72_11_n_1067 & mul_72_11_n_1112)));
 assign mul_72_11_n_1188 = (mul_72_11_n_1098 ^ (mul_72_11_n_1067 ^ mul_72_11_n_1112));
 assign mul_72_11_n_1185 = ((mul_72_11_n_1143 & mul_72_11_n_1101) | ((mul_72_11_n_1101 & mul_72_11_n_1078)
    | (mul_72_11_n_1078 & mul_72_11_n_1143)));
 assign mul_72_11_n_1186 = (mul_72_11_n_1101 ^ (mul_72_11_n_1078 ^ mul_72_11_n_1143));
 assign mul_72_11_n_1183 = ((mul_72_11_n_1099 & mul_72_11_n_1036) | ((mul_72_11_n_1036 & mul_72_11_n_1096)
    | (mul_72_11_n_1096 & mul_72_11_n_1099)));
 assign mul_72_11_n_1184 = (mul_72_11_n_1036 ^ (mul_72_11_n_1096 ^ mul_72_11_n_1099));
 assign mul_72_11_n_1181 = ((mul_72_11_n_1107 & mul_72_11_n_1080) | ((mul_72_11_n_1080 & mul_72_11_n_1090)
    | (mul_72_11_n_1090 & mul_72_11_n_1107)));
 assign mul_72_11_n_1182 = (mul_72_11_n_1080 ^ (mul_72_11_n_1090 ^ mul_72_11_n_1107));
 assign mul_72_11_n_1179 = ((mul_72_11_n_1063 & mul_72_11_n_1126) | ((mul_72_11_n_1126 & mul_72_11_n_1029)
    | (mul_72_11_n_1029 & mul_72_11_n_1063)));
 assign mul_72_11_n_1180 = (mul_72_11_n_1126 ^ (mul_72_11_n_1029 ^ mul_72_11_n_1063));
 assign mul_72_11_n_1177 = ((mul_72_11_n_1109 & mul_72_11_n_1030) | ((mul_72_11_n_1030 & mul_72_11_n_1050)
    | (mul_72_11_n_1050 & mul_72_11_n_1109)));
 assign mul_72_11_n_1178 = (mul_72_11_n_1030 ^ (mul_72_11_n_1050 ^ mul_72_11_n_1109));
 assign mul_72_11_n_1176 = ~(mul_72_11_n_1170 & mul_72_11_n_1173);
 assign mul_72_11_n_1175 = ~(mul_72_11_n_1172 & ~mul_72_11_n_1171);
 assign mul_72_11_n_1174 = ~(mul_72_11_n_1134 | ~mul_72_11_n_1170);
 assign mul_72_11_n_1168 = ((mul_72_11_n_1082 & mul_72_11_n_1083) | ((mul_72_11_n_1083 & mul_72_11_n_995)
    | (mul_72_11_n_995 & mul_72_11_n_1082)));
 assign mul_72_11_n_1169 = (mul_72_11_n_1083 ^ (mul_72_11_n_995 ^ mul_72_11_n_1082));
 assign mul_72_11_n_1166 = ((mul_72_11_n_1092 & mul_72_11_n_1051) | ((mul_72_11_n_1051 & mul_72_11_n_1081)
    | (mul_72_11_n_1081 & mul_72_11_n_1092)));
 assign mul_72_11_n_1167 = (mul_72_11_n_1051 ^ (mul_72_11_n_1081 ^ mul_72_11_n_1092));
 assign mul_72_11_n_1164 = ((mul_72_11_n_1124 & mul_72_11_n_1049) | ((mul_72_11_n_1049 & mul_72_11_n_1037)
    | (mul_72_11_n_1037 & mul_72_11_n_1124)));
 assign mul_72_11_n_1165 = (mul_72_11_n_1049 ^ (mul_72_11_n_1037 ^ mul_72_11_n_1124));
 assign mul_72_11_n_1162 = ((mul_72_11_n_1038 & mul_72_11_n_1077) | ((mul_72_11_n_1077 & mul_72_11_n_1053)
    | (mul_72_11_n_1053 & mul_72_11_n_1038)));
 assign mul_72_11_n_1163 = (mul_72_11_n_1077 ^ (mul_72_11_n_1053 ^ mul_72_11_n_1038));
 assign mul_72_11_n_1173 = ~(mul_72_11_n_1154 & mul_72_11_n_1115);
 assign mul_72_11_n_1172 = ~(mul_72_11_n_1136 & mul_72_11_n_1153);
 assign mul_72_11_n_1171 = ~(mul_72_11_n_1136 | mul_72_11_n_1153);
 assign mul_72_11_n_1170 = (mul_72_11_n_1154 | mul_72_11_n_1115);
 assign {out1[12]} = ~(mul_72_11_n_1145 ^ mul_72_11_n_1089);
 assign mul_72_11_n_1159 = ~(mul_72_11_n_1137 ^ mul_72_11_n_1140);
 assign mul_72_11_n_1158 = ~(mul_72_11_n_1150 & ~mul_72_11_n_1149);
 assign mul_72_11_n_1157 = ~(mul_72_11_n_1073 & (mul_72_11_n_1145 | mul_72_11_n_1075));
 assign mul_72_11_n_1161 = ~(mul_72_11_n_1138 | (mul_72_11_n_1120 & mul_72_11_n_1144));
 assign mul_72_11_n_1155 = ((mul_72_11_n_1065 & mul_72_11_n_1003) | ((mul_72_11_n_1003 & mul_72_11_n_1054)
    | (mul_72_11_n_1054 & mul_72_11_n_1065)));
 assign mul_72_11_n_1156 = (mul_72_11_n_1003 ^ (mul_72_11_n_1054 ^ mul_72_11_n_1065));
 assign mul_72_11_n_1153 = ((mul_72_11_n_1032 & mul_72_11_n_963) | ((mul_72_11_n_963 & mul_72_11_n_1056)
    | (mul_72_11_n_1056 & mul_72_11_n_1032)));
 assign mul_72_11_n_1154 = (mul_72_11_n_963 ^ (mul_72_11_n_1056 ^ mul_72_11_n_1032));
 assign mul_72_11_n_1151 = ((mul_72_11_n_1059 & mul_72_11_n_1091) | ((mul_72_11_n_1091 & mul_72_11_n_1060)
    | (mul_72_11_n_1060 & mul_72_11_n_1059)));
 assign mul_72_11_n_1152 = (mul_72_11_n_1091 ^ (mul_72_11_n_1060 ^ mul_72_11_n_1059));
 assign mul_72_11_n_1150 = ~(mul_72_11_n_1147 & mul_72_11_n_1135);
 assign mul_72_11_n_1149 = ~(mul_72_11_n_1147 | mul_72_11_n_1135);
 assign mul_72_11_n_1148 = ~(mul_72_11_n_1117 ^ mul_72_11_n_1020);
 assign mul_72_11_n_1145 = ~mul_72_11_n_1144;
 assign mul_72_11_n_1142 = ((mul_72_11_n_1028 & mul_72_11_n_1062) | ((mul_72_11_n_1062 & mul_72_11_n_1064)
    | (mul_72_11_n_1064 & mul_72_11_n_1028)));
 assign mul_72_11_n_1143 = (mul_72_11_n_1062 ^ (mul_72_11_n_1064 ^ mul_72_11_n_1028));
 assign mul_72_11_n_1146 = ((mul_72_11_n_1097 & mul_72_11_n_1033) | ((mul_72_11_n_1033 & mul_72_11_n_1001)
    | (mul_72_11_n_1001 & mul_72_11_n_1097)));
 assign mul_72_11_n_1147 = (mul_72_11_n_1033 ^ (mul_72_11_n_1001 ^ mul_72_11_n_1097));
 assign mul_72_11_n_1140 = ((mul_72_11_n_1058 & mul_72_11_n_1024) | ((mul_72_11_n_1024 & mul_72_11_n_998)
    | (mul_72_11_n_998 & mul_72_11_n_1058)));
 assign mul_72_11_n_1141 = (mul_72_11_n_1024 ^ (mul_72_11_n_998 ^ mul_72_11_n_1058));
 assign mul_72_11_n_1139 = ~(mul_72_11_n_1134 | mul_72_11_n_1133);
 assign mul_72_11_n_1144 = ~(mul_72_11_n_1119 & mul_72_11_n_1114);
 assign mul_72_11_n_1138 = ~(mul_72_11_n_1113 & (mul_72_11_n_1106 | mul_72_11_n_1073));
 assign mul_72_11_n_1137 = ~(mul_72_11_n_1105 ^ mul_72_11_n_1008);
 assign mul_72_11_n_1133 = ~mul_72_11_n_1132;
 assign mul_72_11_n_1130 = ((mul_72_11_n_1066 & mul_72_11_n_1016) | ((mul_72_11_n_1016 & mul_72_11_n_1011)
    | (mul_72_11_n_1011 & mul_72_11_n_1066)));
 assign mul_72_11_n_1131 = (mul_72_11_n_1016 ^ (mul_72_11_n_1011 ^ mul_72_11_n_1066));
 assign mul_72_11_n_1128 = ((mul_72_11_n_991 & mul_72_11_n_743) | ((mul_72_11_n_743 & mul_72_11_n_1052)
    | (mul_72_11_n_1052 & mul_72_11_n_991)));
 assign mul_72_11_n_1129 = (mul_72_11_n_743 ^ (mul_72_11_n_1052 ^ mul_72_11_n_991));
 assign mul_72_11_n_1135 = ((mul_72_11_n_1031 & mul_72_11_n_1034) | ((mul_72_11_n_1034 & mul_72_11_n_1015)
    | (mul_72_11_n_1015 & mul_72_11_n_1031)));
 assign mul_72_11_n_1136 = (mul_72_11_n_1034 ^ (mul_72_11_n_1015 ^ mul_72_11_n_1031));
 assign mul_72_11_n_1126 = ((mul_72_11_n_1055 & mul_72_11_n_965) | ((mul_72_11_n_965 & mul_72_11_n_1012)
    | (mul_72_11_n_1012 & mul_72_11_n_1055)));
 assign mul_72_11_n_1127 = (mul_72_11_n_965 ^ (mul_72_11_n_1012 ^ mul_72_11_n_1055));
 assign mul_72_11_n_1124 = ((mul_72_11_n_1027 & mul_72_11_n_735) | ((mul_72_11_n_735 & mul_72_11_n_768)
    | (mul_72_11_n_768 & mul_72_11_n_1027)));
 assign mul_72_11_n_1125 = (mul_72_11_n_735 ^ (mul_72_11_n_768 ^ mul_72_11_n_1027));
 assign mul_72_11_n_1122 = ((mul_72_11_n_1026 & mul_72_11_n_1010) | ((mul_72_11_n_1010 & mul_72_11_n_1046)
    | (mul_72_11_n_1046 & mul_72_11_n_1026)));
 assign mul_72_11_n_1123 = (mul_72_11_n_1010 ^ (mul_72_11_n_1046 ^ mul_72_11_n_1026));
 assign mul_72_11_n_1121 = ~(mul_72_11_n_1113 & ~mul_72_11_n_1106);
 assign mul_72_11_n_1134 = ~(mul_72_11_n_1116 | mul_72_11_n_1103);
 assign mul_72_11_n_1132 = ~(mul_72_11_n_1116 & mul_72_11_n_1103);
 assign {out1[11]} = ~(mul_72_11_n_1085 ^ mul_72_11_n_1088);
 assign mul_72_11_n_1117 = ~(mul_72_11_n_1094 ^ mul_72_11_n_1043);
 assign mul_72_11_n_1120 = ~(mul_72_11_n_1106 | mul_72_11_n_1075);
 assign mul_72_11_n_1119 = ~(mul_72_11_n_1074 | ((mul_72_11_n_1102 & mul_72_11_n_1021) | (mul_72_11_n_1076
    & mul_72_11_n_1040)));
 assign mul_72_11_n_1111 = ((mul_72_11_n_1017 & mul_72_11_n_1035) | ((mul_72_11_n_1035 & mul_72_11_n_945)
    | (mul_72_11_n_945 & mul_72_11_n_1017)));
 assign mul_72_11_n_1112 = (mul_72_11_n_1035 ^ (mul_72_11_n_945 ^ mul_72_11_n_1017));
 assign mul_72_11_n_1115 = ((mul_72_11_n_1057 & mul_72_11_n_952) | ((mul_72_11_n_952 & mul_72_11_n_933)
    | (mul_72_11_n_933 & mul_72_11_n_1057)));
 assign mul_72_11_n_1116 = (mul_72_11_n_952 ^ (mul_72_11_n_933 ^ mul_72_11_n_1057));
 assign mul_72_11_n_1109 = ((mul_72_11_n_1013 & mul_72_11_n_791) | ((mul_72_11_n_791 & mul_72_11_n_994)
    | (mul_72_11_n_994 & mul_72_11_n_1013)));
 assign mul_72_11_n_1110 = (mul_72_11_n_791 ^ (mul_72_11_n_994 ^ mul_72_11_n_1013));
 assign mul_72_11_n_1107 = ((mul_72_11_n_1048 & mul_72_11_n_731) | ((mul_72_11_n_731 & mul_72_11_n_999)
    | (mul_72_11_n_999 & mul_72_11_n_1048)));
 assign mul_72_11_n_1108 = (mul_72_11_n_731 ^ (mul_72_11_n_999 ^ mul_72_11_n_1048));
 assign mul_72_11_n_1114 = ~(mul_72_11_n_1022 & mul_72_11_n_1102);
 assign mul_72_11_n_1113 = ~(mul_72_11_n_1104 & mul_72_11_n_1069);
 assign mul_72_11_n_1105 = ~(mul_72_11_n_1079 ^ mul_72_11_n_1023);
 assign mul_72_11_n_1106 = ~(mul_72_11_n_1104 | mul_72_11_n_1069);
 assign mul_72_11_n_1100 = ((mul_72_11_n_1002 & mul_72_11_n_769) | ((mul_72_11_n_769 & mul_72_11_n_756)
    | (mul_72_11_n_756 & mul_72_11_n_1002)));
 assign mul_72_11_n_1101 = (mul_72_11_n_769 ^ (mul_72_11_n_756 ^ mul_72_11_n_1002));
 assign mul_72_11_n_1098 = ((mul_72_11_n_1000 & mul_72_11_n_982) | ((mul_72_11_n_982 & mul_72_11_n_789)
    | (mul_72_11_n_789 & mul_72_11_n_1000)));
 assign mul_72_11_n_1099 = (mul_72_11_n_982 ^ (mul_72_11_n_789 ^ mul_72_11_n_1000));
 assign mul_72_11_n_1096 = ((mul_72_11_n_939 & mul_72_11_n_737) | ((mul_72_11_n_737 & mul_72_11_n_1014)
    | (mul_72_11_n_1014 & mul_72_11_n_939)));
 assign mul_72_11_n_1097 = (mul_72_11_n_737 ^ (mul_72_11_n_1014 ^ mul_72_11_n_939));
 assign mul_72_11_n_1094 = ((mul_72_11_n_951 & mul_72_11_n_976) | ((mul_72_11_n_976 & mul_72_11_n_915)
    | (mul_72_11_n_915 & mul_72_11_n_951)));
 assign mul_72_11_n_1095 = (mul_72_11_n_976 ^ (mul_72_11_n_915 ^ mul_72_11_n_951));
 assign mul_72_11_n_1103 = ((mul_72_11_n_978 & mul_72_11_n_953) | ((mul_72_11_n_953 & mul_72_11_n_996)
    | (mul_72_11_n_996 & mul_72_11_n_978)));
 assign mul_72_11_n_1104 = (mul_72_11_n_953 ^ (mul_72_11_n_996 ^ mul_72_11_n_978));
 assign mul_72_11_n_1092 = ((mul_72_11_n_1025 & mul_72_11_n_795) | ((mul_72_11_n_795 & mul_72_11_n_751)
    | (mul_72_11_n_751 & mul_72_11_n_1025)));
 assign mul_72_11_n_1093 = (mul_72_11_n_795 ^ (mul_72_11_n_751 ^ mul_72_11_n_1025));
 assign mul_72_11_n_1090 = ((mul_72_11_n_972 & mul_72_11_n_990) | ((mul_72_11_n_990 & mul_72_11_n_742)
    | (mul_72_11_n_742 & mul_72_11_n_972)));
 assign mul_72_11_n_1091 = (mul_72_11_n_990 ^ (mul_72_11_n_742 ^ mul_72_11_n_972));
 assign mul_72_11_n_1089 = ~(mul_72_11_n_1075 | ~mul_72_11_n_1073);
 assign mul_72_11_n_1088 = ~(mul_72_11_n_1076 & ~mul_72_11_n_1074);
 assign mul_72_11_n_1102 = ~(mul_72_11_n_1039 | ~mul_72_11_n_1076);
 assign {out1[10]} = ~(mul_72_11_n_1045 ^ mul_72_11_n_1068);
 assign {out1[9]} = ~(mul_72_11_n_1042 ^ mul_72_11_n_1009);
 assign mul_72_11_n_1085 = ~(mul_72_11_n_1041 & (mul_72_11_n_1068 | mul_72_11_n_1039));
 assign mul_72_11_n_1083 = ((mul_72_11_n_974 & mul_72_11_n_796) | ((mul_72_11_n_796 & mul_72_11_n_772)
    | (mul_72_11_n_772 & mul_72_11_n_974)));
 assign mul_72_11_n_1084 = (mul_72_11_n_796 ^ (mul_72_11_n_772 ^ mul_72_11_n_974));
 assign mul_72_11_n_1081 = ((mul_72_11_n_973 & mul_72_11_n_955) | ((mul_72_11_n_955 & mul_72_11_n_916)
    | (mul_72_11_n_916 & mul_72_11_n_973)));
 assign mul_72_11_n_1082 = (mul_72_11_n_955 ^ (mul_72_11_n_916 ^ mul_72_11_n_973));
 assign mul_72_11_n_1079 = ((mul_72_11_n_971 & mul_72_11_n_730) | ((mul_72_11_n_730 & mul_72_11_n_763)
    | (mul_72_11_n_763 & mul_72_11_n_971)));
 assign mul_72_11_n_1080 = (mul_72_11_n_730 ^ (mul_72_11_n_763 ^ mul_72_11_n_971));
 assign mul_72_11_n_1077 = ((mul_72_11_n_993 & mul_72_11_n_759) | ((mul_72_11_n_759 & mul_72_11_n_946)
    | (mul_72_11_n_946 & mul_72_11_n_993)));
 assign mul_72_11_n_1078 = (mul_72_11_n_759 ^ (mul_72_11_n_946 ^ mul_72_11_n_993));
 assign mul_72_11_n_1076 = (mul_72_11_n_1072 | mul_72_11_n_1018);
 assign mul_72_11_n_1075 = ~(mul_72_11_n_1070 | mul_72_11_n_1071);
 assign mul_72_11_n_1074 = (mul_72_11_n_1072 & mul_72_11_n_1018);
 assign mul_72_11_n_1073 = ~(mul_72_11_n_1070 & mul_72_11_n_1071);
 assign mul_72_11_n_1066 = ((mul_72_11_n_913 & mul_72_11_n_981) | ((mul_72_11_n_981 & mul_72_11_n_788)
    | (mul_72_11_n_788 & mul_72_11_n_913)));
 assign mul_72_11_n_1067 = (mul_72_11_n_981 ^ (mul_72_11_n_788 ^ mul_72_11_n_913));
 assign mul_72_11_n_1064 = ((mul_72_11_n_908 & mul_72_11_n_947) | ((mul_72_11_n_947 & mul_72_11_n_979)
    | (mul_72_11_n_979 & mul_72_11_n_908)));
 assign mul_72_11_n_1065 = (mul_72_11_n_947 ^ (mul_72_11_n_979 ^ mul_72_11_n_908));
 assign mul_72_11_n_1062 = ((mul_72_11_n_961 & mul_72_11_n_757) | ((mul_72_11_n_757 & mul_72_11_n_964)
    | (mul_72_11_n_964 & mul_72_11_n_961)));
 assign mul_72_11_n_1063 = (mul_72_11_n_757 ^ (mul_72_11_n_964 ^ mul_72_11_n_961));
 assign mul_72_11_n_1060 = ((mul_72_11_n_957 & mul_72_11_n_734) | ((mul_72_11_n_734 & mul_72_11_n_744)
    | (mul_72_11_n_744 & mul_72_11_n_957)));
 assign mul_72_11_n_1061 = (mul_72_11_n_734 ^ (mul_72_11_n_744 ^ mul_72_11_n_957));
 assign mul_72_11_n_1058 = ((mul_72_11_n_923 & mul_72_11_n_927) | ((mul_72_11_n_927 & mul_72_11_n_956)
    | (mul_72_11_n_956 & mul_72_11_n_923)));
 assign mul_72_11_n_1059 = (mul_72_11_n_927 ^ (mul_72_11_n_956 ^ mul_72_11_n_923));
 assign mul_72_11_n_1056 = ((mul_72_11_n_893 & mul_72_11_n_888) | ((mul_72_11_n_888 & mul_72_11_n_977)
    | (mul_72_11_n_977 & mul_72_11_n_893)));
 assign mul_72_11_n_1057 = (mul_72_11_n_888 ^ (mul_72_11_n_977 ^ mul_72_11_n_893));
 assign mul_72_11_n_1054 = ((mul_72_11_n_958 & mul_72_11_n_930) | ((mul_72_11_n_930 & mul_72_11_n_660)
    | (mul_72_11_n_660 & mul_72_11_n_958)));
 assign mul_72_11_n_1055 = (mul_72_11_n_930 ^ (mul_72_11_n_660 ^ mul_72_11_n_958));
 assign mul_72_11_n_1052 = ((mul_72_11_n_992 & mul_72_11_n_758) | ((mul_72_11_n_758 & mul_72_11_n_904)
    | (mul_72_11_n_904 & mul_72_11_n_992)));
 assign mul_72_11_n_1053 = (mul_72_11_n_758 ^ (mul_72_11_n_904 ^ mul_72_11_n_992));
 assign mul_72_11_n_1050 = ((mul_72_11_n_959 & mul_72_11_n_931) | ((mul_72_11_n_931 & mul_72_11_n_750)
    | (mul_72_11_n_750 & mul_72_11_n_959)));
 assign mul_72_11_n_1051 = (mul_72_11_n_931 ^ (mul_72_11_n_750 ^ mul_72_11_n_959));
 assign mul_72_11_n_1071 = ((mul_72_11_n_921 & mul_72_11_n_924) | ((mul_72_11_n_924 & mul_72_11_n_883)
    | (mul_72_11_n_883 & mul_72_11_n_921)));
 assign mul_72_11_n_1072 = (mul_72_11_n_924 ^ (mul_72_11_n_883 ^ mul_72_11_n_921));
 assign mul_72_11_n_1048 = ((mul_72_11_n_918 & mul_72_11_n_771) | ((mul_72_11_n_771 & mul_72_11_n_928)
    | (mul_72_11_n_928 & mul_72_11_n_918)));
 assign mul_72_11_n_1049 = (mul_72_11_n_771 ^ (mul_72_11_n_928 ^ mul_72_11_n_918));
 assign mul_72_11_n_1069 = ((mul_72_11_n_997 & mul_72_11_n_733) | ((mul_72_11_n_733 & mul_72_11_n_920)
    | (mul_72_11_n_920 & mul_72_11_n_997)));
 assign mul_72_11_n_1070 = (mul_72_11_n_733 ^ (mul_72_11_n_920 ^ mul_72_11_n_997));
 assign mul_72_11_n_1046 = ((mul_72_11_n_949 & mul_72_11_n_773) | ((mul_72_11_n_773 & mul_72_11_n_944)
    | (mul_72_11_n_944 & mul_72_11_n_949)));
 assign mul_72_11_n_1047 = (mul_72_11_n_773 ^ (mul_72_11_n_944 ^ mul_72_11_n_949));
 assign mul_72_11_n_1045 = ~(mul_72_11_n_1039 | mul_72_11_n_1040);
 assign mul_72_11_n_1068 = ~(mul_72_11_n_1022 | mul_72_11_n_1021);
 assign {out1[8]} = ~(mul_72_11_n_1007 ^ mul_72_11_n_989);
 assign mul_72_11_n_1043 = ~(mul_72_11_n_1006 ^ mul_72_11_n_910);
 assign mul_72_11_n_1042 = ~(mul_72_11_n_983 & (mul_72_11_n_1007 | mul_72_11_n_970));
 assign mul_72_11_n_1041 = ~mul_72_11_n_1040;
 assign mul_72_11_n_1037 = ((mul_72_11_n_929 & mul_72_11_n_745) | ((mul_72_11_n_745 & mul_72_11_n_919)
    | (mul_72_11_n_919 & mul_72_11_n_929)));
 assign mul_72_11_n_1038 = (mul_72_11_n_745 ^ (mul_72_11_n_919 ^ mul_72_11_n_929));
 assign mul_72_11_n_1035 = ((mul_72_11_n_938 & mul_72_11_n_736) | ((mul_72_11_n_736 & mul_72_11_n_901)
    | (mul_72_11_n_901 & mul_72_11_n_938)));
 assign mul_72_11_n_1036 = (mul_72_11_n_736 ^ (mul_72_11_n_901 ^ mul_72_11_n_938));
 assign mul_72_11_n_1033 = ((mul_72_11_n_937 & mul_72_11_n_962) | ((mul_72_11_n_962 & mul_72_11_n_934)
    | (mul_72_11_n_934 & mul_72_11_n_937)));
 assign mul_72_11_n_1034 = (mul_72_11_n_962 ^ (mul_72_11_n_934 ^ mul_72_11_n_937));
 assign mul_72_11_n_1031 = ((mul_72_11_n_935 & mul_72_11_n_932) | ((mul_72_11_n_932 & mul_72_11_n_895)
    | (mul_72_11_n_895 & mul_72_11_n_935)));
 assign mul_72_11_n_1032 = (mul_72_11_n_932 ^ (mul_72_11_n_895 ^ mul_72_11_n_935));
 assign mul_72_11_n_1029 = ((mul_72_11_n_980 & mul_72_11_n_790) | ((mul_72_11_n_790 & mul_72_11_n_909)
    | (mul_72_11_n_909 & mul_72_11_n_980)));
 assign mul_72_11_n_1030 = (mul_72_11_n_790 ^ (mul_72_11_n_909 ^ mul_72_11_n_980));
 assign mul_72_11_n_1027 = ((mul_72_11_n_905 & mul_72_11_n_519) | ((mul_72_11_n_519 & mul_72_11_n_960)
    | (mul_72_11_n_960 & mul_72_11_n_905)));
 assign mul_72_11_n_1028 = (mul_72_11_n_519 ^ (mul_72_11_n_960 ^ mul_72_11_n_905));
 assign mul_72_11_n_1025 = ((mul_72_11_n_917 & mul_72_11_n_948) | ((mul_72_11_n_948 & mul_72_11_n_511)
    | (mul_72_11_n_511 & mul_72_11_n_917)));
 assign mul_72_11_n_1026 = (mul_72_11_n_948 ^ (mul_72_11_n_511 ^ mul_72_11_n_917));
 assign mul_72_11_n_1023 = ((mul_72_11_n_922 & mul_72_11_n_926) | ((mul_72_11_n_926 & mul_72_11_n_663)
    | (mul_72_11_n_663 & mul_72_11_n_922)));
 assign mul_72_11_n_1024 = (mul_72_11_n_926 ^ (mul_72_11_n_663 ^ mul_72_11_n_922));
 assign mul_72_11_n_1040 = (mul_72_11_n_1019 & mul_72_11_n_984);
 assign mul_72_11_n_1039 = ~(mul_72_11_n_1019 | mul_72_11_n_984);
 assign mul_72_11_n_1022 = ~(mul_72_11_n_1004 | (mul_72_11_n_970 | mul_72_11_n_1007));
 assign mul_72_11_n_1021 = ~(mul_72_11_n_1005 & (mul_72_11_n_1004 | mul_72_11_n_983));
 assign mul_72_11_n_1020 = ~(mul_72_11_n_986 ^ mul_72_11_n_727);
 assign mul_72_11_n_1016 = ((mul_72_11_n_900 & mul_72_11_n_497) | ((mul_72_11_n_497 & mul_72_11_n_897)
    | (mul_72_11_n_897 & mul_72_11_n_900)));
 assign mul_72_11_n_1017 = (mul_72_11_n_497 ^ (mul_72_11_n_897 ^ mul_72_11_n_900));
 assign mul_72_11_n_1014 = ((mul_72_11_n_867 & mul_72_11_n_894) | ((mul_72_11_n_894 & mul_72_11_n_827)
    | (mul_72_11_n_827 & mul_72_11_n_867)));
 assign mul_72_11_n_1015 = (mul_72_11_n_894 ^ (mul_72_11_n_827 ^ mul_72_11_n_867));
 assign mul_72_11_n_1018 = ((mul_72_11_n_925 & mul_72_11_n_886) | ((mul_72_11_n_886 & mul_72_11_n_844)
    | (mul_72_11_n_844 & mul_72_11_n_925)));
 assign mul_72_11_n_1019 = (mul_72_11_n_886 ^ (mul_72_11_n_844 ^ mul_72_11_n_925));
 assign mul_72_11_n_1012 = ((mul_72_11_n_954 & mul_72_11_n_884) | ((mul_72_11_n_884 & mul_72_11_n_507)
    | (mul_72_11_n_507 & mul_72_11_n_954)));
 assign mul_72_11_n_1013 = (mul_72_11_n_884 ^ (mul_72_11_n_507 ^ mul_72_11_n_954));
 assign mul_72_11_n_1010 = ((mul_72_11_n_912 & mul_72_11_n_729) | ((mul_72_11_n_729 & mul_72_11_n_896)
    | (mul_72_11_n_896 & mul_72_11_n_912)));
 assign mul_72_11_n_1011 = (mul_72_11_n_729 ^ (mul_72_11_n_896 ^ mul_72_11_n_912));
 assign mul_72_11_n_1009 = ~(mul_72_11_n_1005 & ~mul_72_11_n_1004);
 assign mul_72_11_n_1008 = ~(mul_72_11_n_969 ^ mul_72_11_n_855);
 assign mul_72_11_n_1006 = ~(mul_72_11_n_975 ^ mul_72_11_n_875);
 assign mul_72_11_n_1007 = ~(mul_72_11_n_988 | ((mul_72_11_n_911 & mul_72_11_n_857) | (mul_72_11_n_966
    & mul_72_11_n_874)));
 assign mul_72_11_n_1002 = ((mul_72_11_n_898 & mul_72_11_n_661) | ((mul_72_11_n_661 & mul_72_11_n_516)
    | (mul_72_11_n_516 & mul_72_11_n_898)));
 assign mul_72_11_n_1003 = (mul_72_11_n_661 ^ (mul_72_11_n_516 ^ mul_72_11_n_898));
 assign mul_72_11_n_1000 = ((mul_72_11_n_936 & mul_72_11_n_866) | ((mul_72_11_n_866 & mul_72_11_n_873)
    | (mul_72_11_n_873 & mul_72_11_n_936)));
 assign mul_72_11_n_1001 = (mul_72_11_n_866 ^ (mul_72_11_n_873 ^ mul_72_11_n_936));
 assign mul_72_11_n_998 = ((mul_72_11_n_890 & mul_72_11_n_770) | ((mul_72_11_n_770 & mul_72_11_n_668)
    | (mul_72_11_n_668 & mul_72_11_n_890)));
 assign mul_72_11_n_999 = (mul_72_11_n_770 ^ (mul_72_11_n_668 ^ mul_72_11_n_890));
 assign mul_72_11_n_996 = ((mul_72_11_n_882 & mul_72_11_n_807) | ((mul_72_11_n_807 & mul_72_11_n_842)
    | (mul_72_11_n_842 & mul_72_11_n_882)));
 assign mul_72_11_n_997 = (mul_72_11_n_807 ^ (mul_72_11_n_842 ^ mul_72_11_n_882));
 assign mul_72_11_n_994 = ((mul_72_11_n_885 & mul_72_11_n_506) | ((mul_72_11_n_506 & mul_72_11_n_862)
    | (mul_72_11_n_862 & mul_72_11_n_885)));
 assign mul_72_11_n_995 = (mul_72_11_n_506 ^ (mul_72_11_n_862 ^ mul_72_11_n_885));
 assign mul_72_11_n_992 = ((mul_72_11_n_829 & mul_72_11_n_503) | ((mul_72_11_n_503 & mul_72_11_n_878)
    | (mul_72_11_n_878 & mul_72_11_n_829)));
 assign mul_72_11_n_993 = (mul_72_11_n_503 ^ (mul_72_11_n_878 ^ mul_72_11_n_829));
 assign mul_72_11_n_990 = ((mul_72_11_n_891 & mul_72_11_n_662) | ((mul_72_11_n_662 & mul_72_11_n_638)
    | (mul_72_11_n_638 & mul_72_11_n_891)));
 assign mul_72_11_n_991 = (mul_72_11_n_662 ^ (mul_72_11_n_638 ^ mul_72_11_n_891));
 assign mul_72_11_n_989 = ~(mul_72_11_n_970 | ~mul_72_11_n_983);
 assign mul_72_11_n_1005 = ~(mul_72_11_n_985 & mul_72_11_n_967);
 assign mul_72_11_n_1004 = ~(mul_72_11_n_985 | mul_72_11_n_967);
 assign mul_72_11_n_988 = ~(mul_72_11_n_940 & ~(mul_72_11_n_966 & mul_72_11_n_876));
 assign {out1[7]} = ~(mul_72_11_n_943 ^ mul_72_11_n_941);
 assign mul_72_11_n_986 = ~(mul_72_11_n_697 ^ mul_72_11_n_950);
 assign mul_72_11_n_981 = ((mul_72_11_n_840 & mul_72_11_n_650) | ((mul_72_11_n_650 & mul_72_11_n_872)
    | (mul_72_11_n_872 & mul_72_11_n_840)));
 assign mul_72_11_n_982 = (mul_72_11_n_650 ^ (mul_72_11_n_872 ^ mul_72_11_n_840));
 assign mul_72_11_n_979 = ((mul_72_11_n_868 & mul_72_11_n_646) | ((mul_72_11_n_646 & mul_72_11_n_382)
    | (mul_72_11_n_382 & mul_72_11_n_868)));
 assign mul_72_11_n_980 = (mul_72_11_n_646 ^ (mul_72_11_n_382 ^ mul_72_11_n_868));
 assign mul_72_11_n_977 = ((mul_72_11_n_815 & mul_72_11_n_473) | ((mul_72_11_n_473 & mul_72_11_n_841)
    | (mul_72_11_n_841 & mul_72_11_n_815)));
 assign mul_72_11_n_978 = (mul_72_11_n_473 ^ (mul_72_11_n_841 ^ mul_72_11_n_815));
 assign mul_72_11_n_984 = ((mul_72_11_n_887 & mul_72_11_n_845) | ((mul_72_11_n_845 & mul_72_11_n_825)
    | (mul_72_11_n_825 & mul_72_11_n_887)));
 assign mul_72_11_n_985 = (mul_72_11_n_845 ^ (mul_72_11_n_825 ^ mul_72_11_n_887));
 assign mul_72_11_n_975 = ((mul_72_11_n_864 & mul_72_11_n_514) | ((mul_72_11_n_514 & mul_72_11_n_522)
    | (mul_72_11_n_522 & mul_72_11_n_864)));
 assign mul_72_11_n_976 = (mul_72_11_n_514 ^ (mul_72_11_n_522 ^ mul_72_11_n_864));
 assign mul_72_11_n_973 = ((mul_72_11_n_863 & mul_72_11_n_641) | ((mul_72_11_n_641 & mul_72_11_n_837)
    | (mul_72_11_n_837 & mul_72_11_n_863)));
 assign mul_72_11_n_974 = (mul_72_11_n_641 ^ (mul_72_11_n_837 ^ mul_72_11_n_863));
 assign mul_72_11_n_971 = ((mul_72_11_n_865 & mul_72_11_n_637) | ((mul_72_11_n_637 & mul_72_11_n_647)
    | (mul_72_11_n_647 & mul_72_11_n_865)));
 assign mul_72_11_n_972 = (mul_72_11_n_637 ^ (mul_72_11_n_647 ^ mul_72_11_n_865));
 assign mul_72_11_n_983 = ~(mul_72_11_n_968 & mul_72_11_n_906);
 assign mul_72_11_n_969 = ~(mul_72_11_n_914 ^ mul_72_11_n_762);
 assign mul_72_11_n_970 = ~(mul_72_11_n_968 | mul_72_11_n_906);
 assign mul_72_11_n_964 = ((mul_72_11_n_899 & mul_72_11_n_512) | ((mul_72_11_n_512 & mul_72_11_n_495)
    | (mul_72_11_n_495 & mul_72_11_n_899)));
 assign mul_72_11_n_965 = (mul_72_11_n_512 ^ (mul_72_11_n_495 ^ mul_72_11_n_899));
 assign mul_72_11_n_962 = ((mul_72_11_n_892 & mul_72_11_n_631) | ((mul_72_11_n_631 & mul_72_11_n_578)
    | (mul_72_11_n_578 & mul_72_11_n_892)));
 assign mul_72_11_n_963 = (mul_72_11_n_631 ^ (mul_72_11_n_578 ^ mul_72_11_n_892));
 assign mul_72_11_n_960 = ((mul_72_11_n_806 & mul_72_11_n_849) | ((mul_72_11_n_849 & mul_72_11_n_585)
    | (mul_72_11_n_585 & mul_72_11_n_806)));
 assign mul_72_11_n_961 = (mul_72_11_n_849 ^ (mul_72_11_n_585 ^ mul_72_11_n_806));
 assign mul_72_11_n_958 = ((mul_72_11_n_847 & mul_72_11_n_629) | ((mul_72_11_n_629 & mul_72_11_n_869)
    | (mul_72_11_n_869 & mul_72_11_n_847)));
 assign mul_72_11_n_959 = (mul_72_11_n_629 ^ (mul_72_11_n_869 ^ mul_72_11_n_847));
 assign mul_72_11_n_956 = ((mul_72_11_n_800 & mul_72_11_n_655) | ((mul_72_11_n_655 & mul_72_11_n_870)
    | (mul_72_11_n_870 & mul_72_11_n_800)));
 assign mul_72_11_n_957 = (mul_72_11_n_655 ^ (mul_72_11_n_870 ^ mul_72_11_n_800));
 assign mul_72_11_n_954 = ((mul_72_11_n_848 & mul_72_11_n_400) | ((mul_72_11_n_400 & mul_72_11_n_643)
    | (mul_72_11_n_643 & mul_72_11_n_848)));
 assign mul_72_11_n_955 = (mul_72_11_n_400 ^ (mul_72_11_n_643 ^ mul_72_11_n_848));
 assign mul_72_11_n_967 = ((mul_72_11_n_846 & mul_72_11_n_810) | ((mul_72_11_n_810 & mul_72_11_n_586)
    | (mul_72_11_n_586 & mul_72_11_n_846)));
 assign mul_72_11_n_968 = (mul_72_11_n_810 ^ (mul_72_11_n_586 ^ mul_72_11_n_846));
 assign mul_72_11_n_952 = ((mul_72_11_n_889 & mul_72_11_n_570) | ((mul_72_11_n_570 & mul_72_11_n_732)
    | (mul_72_11_n_732 & mul_72_11_n_889)));
 assign mul_72_11_n_953 = (mul_72_11_n_570 ^ (mul_72_11_n_732 ^ mul_72_11_n_889));
 assign mul_72_11_n_950 = ((mul_72_11_n_881 & mul_72_11_n_667) | ((mul_72_11_n_667 & mul_72_11_n_635)
    | (mul_72_11_n_635 & mul_72_11_n_881)));
 assign mul_72_11_n_951 = (mul_72_11_n_667 ^ (mul_72_11_n_635 ^ mul_72_11_n_881));
 assign mul_72_11_n_948 = ((mul_72_11_n_838 & mul_72_11_n_623) | ((mul_72_11_n_623 & mul_72_11_n_801)
    | (mul_72_11_n_801 & mul_72_11_n_838)));
 assign mul_72_11_n_949 = (mul_72_11_n_623 ^ (mul_72_11_n_801 ^ mul_72_11_n_838));
 assign mul_72_11_n_946 = ((mul_72_11_n_879 & mul_72_11_n_559) | ((mul_72_11_n_559 & mul_72_11_n_633)
    | (mul_72_11_n_633 & mul_72_11_n_879)));
 assign mul_72_11_n_947 = (mul_72_11_n_559 ^ (mul_72_11_n_633 ^ mul_72_11_n_879));
 assign mul_72_11_n_944 = ((mul_72_11_n_839 & mul_72_11_n_652) | ((mul_72_11_n_652 & mul_72_11_n_639)
    | (mul_72_11_n_639 & mul_72_11_n_839)));
 assign mul_72_11_n_945 = (mul_72_11_n_652 ^ (mul_72_11_n_639 ^ mul_72_11_n_839));
 assign mul_72_11_n_943 = ~(mul_72_11_n_911 & mul_72_11_n_940);
 assign mul_72_11_n_966 = ~(mul_72_11_n_859 | ~mul_72_11_n_911);
 assign {out1[6]} = ~(mul_72_11_n_903 ^ mul_72_11_n_877);
 assign mul_72_11_n_941 = ~(mul_72_11_n_858 & (mul_72_11_n_903 | mul_72_11_n_859));
 assign mul_72_11_n_938 = ((mul_72_11_n_831 & mul_72_11_n_480) | ((mul_72_11_n_480 & mul_72_11_n_826)
    | (mul_72_11_n_826 & mul_72_11_n_831)));
 assign mul_72_11_n_939 = (mul_72_11_n_480 ^ (mul_72_11_n_826 ^ mul_72_11_n_831));
 assign mul_72_11_n_936 = ((mul_72_11_n_816 & mul_72_11_n_632) | ((mul_72_11_n_632 & mul_72_11_n_581)
    | (mul_72_11_n_581 & mul_72_11_n_816)));
 assign mul_72_11_n_937 = (mul_72_11_n_632 ^ (mul_72_11_n_581 ^ mul_72_11_n_816));
 assign mul_72_11_n_934 = ((mul_72_11_n_817 & mul_72_11_n_818) | ((mul_72_11_n_818 & mul_72_11_n_476)
    | (mul_72_11_n_476 & mul_72_11_n_817)));
 assign mul_72_11_n_935 = (mul_72_11_n_818 ^ (mul_72_11_n_476 ^ mul_72_11_n_817));
 assign mul_72_11_n_932 = ((mul_72_11_n_819 & mul_72_11_n_625) | ((mul_72_11_n_625 & mul_72_11_n_814)
    | (mul_72_11_n_814 & mul_72_11_n_819)));
 assign mul_72_11_n_933 = (mul_72_11_n_625 ^ (mul_72_11_n_814 ^ mul_72_11_n_819));
 assign mul_72_11_n_930 = ((mul_72_11_n_798 & mul_72_11_n_665) | ((mul_72_11_n_665 & mul_72_11_n_574)
    | (mul_72_11_n_574 & mul_72_11_n_798)));
 assign mul_72_11_n_931 = (mul_72_11_n_665 ^ (mul_72_11_n_574 ^ mul_72_11_n_798));
 assign mul_72_11_n_928 = ((mul_72_11_n_823 & mul_72_11_n_569) | ((mul_72_11_n_569 & mul_72_11_n_828)
    | (mul_72_11_n_828 & mul_72_11_n_823)));
 assign mul_72_11_n_929 = (mul_72_11_n_569 ^ (mul_72_11_n_828 ^ mul_72_11_n_823));
 assign mul_72_11_n_926 = ((mul_72_11_n_799 & mul_72_11_n_492) | ((mul_72_11_n_492 & mul_72_11_n_644)
    | (mul_72_11_n_644 & mul_72_11_n_799)));
 assign mul_72_11_n_927 = (mul_72_11_n_492 ^ (mul_72_11_n_644 ^ mul_72_11_n_799));
 assign mul_72_11_n_924 = ((mul_72_11_n_824 & mul_72_11_n_451) | ((mul_72_11_n_451 & mul_72_11_n_590)
    | (mul_72_11_n_590 & mul_72_11_n_824)));
 assign mul_72_11_n_925 = (mul_72_11_n_451 ^ (mul_72_11_n_590 ^ mul_72_11_n_824));
 assign mul_72_11_n_922 = ((mul_72_11_n_821 & mul_72_11_n_654) | ((mul_72_11_n_654 & mul_72_11_n_576)
    | (mul_72_11_n_576 & mul_72_11_n_821)));
 assign mul_72_11_n_923 = (mul_72_11_n_654 ^ (mul_72_11_n_576 ^ mul_72_11_n_821));
 assign mul_72_11_n_920 = ((mul_72_11_n_808 & mul_72_11_n_843) | ((mul_72_11_n_843 & mul_72_11_n_440)
    | (mul_72_11_n_440 & mul_72_11_n_808)));
 assign mul_72_11_n_921 = (mul_72_11_n_843 ^ (mul_72_11_n_440 ^ mul_72_11_n_808));
 assign mul_72_11_n_918 = ((mul_72_11_n_871 & mul_72_11_n_669) | ((mul_72_11_n_669 & mul_72_11_n_640)
    | (mul_72_11_n_640 & mul_72_11_n_871)));
 assign mul_72_11_n_919 = (mul_72_11_n_669 ^ (mul_72_11_n_640 ^ mul_72_11_n_871));
 assign mul_72_11_n_916 = ((mul_72_11_n_813 & mul_72_11_n_558) | ((mul_72_11_n_558 & mul_72_11_n_624)
    | (mul_72_11_n_624 & mul_72_11_n_813)));
 assign mul_72_11_n_917 = (mul_72_11_n_558 ^ (mul_72_11_n_624 ^ mul_72_11_n_813));
 assign mul_72_11_n_914 = ((mul_72_11_n_804 & mul_72_11_n_502) | ((mul_72_11_n_502 & mul_72_11_n_657)
    | (mul_72_11_n_657 & mul_72_11_n_804)));
 assign mul_72_11_n_915 = (mul_72_11_n_502 ^ (mul_72_11_n_657 ^ mul_72_11_n_804));
 assign mul_72_11_n_912 = ((mul_72_11_n_802 & mul_72_11_n_557) | ((mul_72_11_n_557 & mul_72_11_n_575)
    | (mul_72_11_n_575 & mul_72_11_n_802)));
 assign mul_72_11_n_913 = (mul_72_11_n_557 ^ (mul_72_11_n_575 ^ mul_72_11_n_802));
 assign mul_72_11_n_940 = ~(mul_72_11_n_907 & mul_72_11_n_853);
 assign mul_72_11_n_910 = ~(mul_72_11_n_694 ^ mul_72_11_n_880);
 assign mul_72_11_n_911 = (mul_72_11_n_907 | mul_72_11_n_853);
 assign mul_72_11_n_908 = ((mul_72_11_n_850 & mul_72_11_n_628) | ((mul_72_11_n_628 & mul_72_11_n_577)
    | (mul_72_11_n_577 & mul_72_11_n_850)));
 assign mul_72_11_n_909 = (mul_72_11_n_628 ^ (mul_72_11_n_577 ^ mul_72_11_n_850));
 assign mul_72_11_n_906 = ((mul_72_11_n_811 & mul_72_11_n_567) | ((mul_72_11_n_567 & mul_72_11_n_786)
    | (mul_72_11_n_786 & mul_72_11_n_811)));
 assign mul_72_11_n_907 = (mul_72_11_n_567 ^ (mul_72_11_n_786 ^ mul_72_11_n_811));
 assign mul_72_11_n_904 = ((mul_72_11_n_749 & mul_72_11_n_455) | ((mul_72_11_n_455 & mul_72_11_n_805)
    | (mul_72_11_n_805 & mul_72_11_n_749)));
 assign mul_72_11_n_905 = (mul_72_11_n_455 ^ (mul_72_11_n_805 ^ mul_72_11_n_749));
 assign mul_72_11_n_903 = ~(mul_72_11_n_876 | mul_72_11_n_874);
 assign {out1[5]} = ~(mul_72_11_n_861 ^ mul_72_11_n_860);
 assign mul_72_11_n_900 = ((mul_72_11_n_830 & mul_72_11_n_481) | ((mul_72_11_n_481 & mul_72_11_n_461)
    | (mul_72_11_n_461 & mul_72_11_n_830)));
 assign mul_72_11_n_901 = (mul_72_11_n_481 ^ (mul_72_11_n_461 ^ mul_72_11_n_830));
 assign mul_72_11_n_898 = ((mul_72_11_n_797 & mul_72_11_n_477) | ((mul_72_11_n_477 & mul_72_11_n_449)
    | (mul_72_11_n_449 & mul_72_11_n_797)));
 assign mul_72_11_n_899 = (mul_72_11_n_477 ^ (mul_72_11_n_449 ^ mul_72_11_n_797));
 assign mul_72_11_n_896 = ((mul_72_11_n_774 & mul_72_11_n_435) | ((mul_72_11_n_435 & mul_72_11_n_463)
    | (mul_72_11_n_463 & mul_72_11_n_774)));
 assign mul_72_11_n_897 = (mul_72_11_n_435 ^ (mul_72_11_n_463 ^ mul_72_11_n_774));
 assign mul_72_11_n_894 = ((mul_72_11_n_782 & mul_72_11_n_672) | ((mul_72_11_n_672 & mul_72_11_n_456)
    | (mul_72_11_n_456 & mul_72_11_n_782)));
 assign mul_72_11_n_895 = (mul_72_11_n_672 ^ (mul_72_11_n_456 ^ mul_72_11_n_782));
 assign mul_72_11_n_892 = ((mul_72_11_n_783 & mul_72_11_n_403) | ((mul_72_11_n_403 & mul_72_11_n_478)
    | (mul_72_11_n_478 & mul_72_11_n_783)));
 assign mul_72_11_n_893 = (mul_72_11_n_403 ^ (mul_72_11_n_478 ^ mul_72_11_n_783));
 assign mul_72_11_n_890 = ((mul_72_11_n_822 & mul_72_11_n_472) | ((mul_72_11_n_472 & mul_72_11_n_741)
    | (mul_72_11_n_741 & mul_72_11_n_822)));
 assign mul_72_11_n_891 = (mul_72_11_n_472 ^ (mul_72_11_n_741 ^ mul_72_11_n_822));
 assign mul_72_11_n_888 = ((mul_72_11_n_784 & mul_72_11_n_671) | ((mul_72_11_n_671 & mul_72_11_n_454)
    | (mul_72_11_n_454 & mul_72_11_n_784)));
 assign mul_72_11_n_889 = (mul_72_11_n_671 ^ (mul_72_11_n_454 ^ mul_72_11_n_784));
 assign mul_72_11_n_886 = ((mul_72_11_n_776 & mul_72_11_n_452) | ((mul_72_11_n_452 & mul_72_11_n_591)
    | (mul_72_11_n_591 & mul_72_11_n_776)));
 assign mul_72_11_n_887 = (mul_72_11_n_452 ^ (mul_72_11_n_591 ^ mul_72_11_n_776));
 assign mul_72_11_n_884 = ((mul_72_11_n_812 & mul_72_11_n_470) | ((mul_72_11_n_470 & mul_72_11_n_448)
    | (mul_72_11_n_448 & mul_72_11_n_812)));
 assign mul_72_11_n_885 = (mul_72_11_n_470 ^ (mul_72_11_n_448 ^ mul_72_11_n_812));
 assign mul_72_11_n_882 = ((mul_72_11_n_778 & mul_72_11_n_447) | ((mul_72_11_n_447 & mul_72_11_n_589)
    | (mul_72_11_n_589 & mul_72_11_n_778)));
 assign mul_72_11_n_883 = (mul_72_11_n_447 ^ (mul_72_11_n_589 ^ mul_72_11_n_778));
 assign mul_72_11_n_880 = ((mul_72_11_n_820 & mul_72_11_n_491) | ((mul_72_11_n_491 & mul_72_11_n_739)
    | (mul_72_11_n_739 & mul_72_11_n_820)));
 assign mul_72_11_n_881 = (mul_72_11_n_491 ^ (mul_72_11_n_739 ^ mul_72_11_n_820));
 assign mul_72_11_n_878 = ((mul_72_11_n_780 & mul_72_11_n_457) | ((mul_72_11_n_457 & mul_72_11_n_464)
    | (mul_72_11_n_464 & mul_72_11_n_780)));
 assign mul_72_11_n_879 = (mul_72_11_n_457 ^ (mul_72_11_n_464 ^ mul_72_11_n_780));
 assign mul_72_11_n_877 = ~(mul_72_11_n_859 | mul_72_11_n_857);
 assign mul_72_11_n_876 = ~(mul_72_11_n_852 & (mul_72_11_n_851 | mul_72_11_n_767));
 assign mul_72_11_n_875 = ~(mul_72_11_n_766 ^ mul_72_11_n_835);
 assign mul_72_11_n_872 = ((mul_72_11_n_754 & mul_72_11_n_653) | ((mul_72_11_n_653 & mul_72_11_n_460)
    | (mul_72_11_n_460 & mul_72_11_n_754)));
 assign mul_72_11_n_873 = (mul_72_11_n_653 ^ (mul_72_11_n_460 ^ mul_72_11_n_754));
 assign mul_72_11_n_870 = ((mul_72_11_n_748 & mul_72_11_n_465) | ((mul_72_11_n_465 & mul_72_11_n_468)
    | (mul_72_11_n_468 & mul_72_11_n_748)));
 assign mul_72_11_n_871 = (mul_72_11_n_465 ^ (mul_72_11_n_468 ^ mul_72_11_n_748));
 assign mul_72_11_n_868 = ((mul_72_11_n_752 & mul_72_11_n_475) | ((mul_72_11_n_475 & mul_72_11_n_434)
    | (mul_72_11_n_434 & mul_72_11_n_752)));
 assign mul_72_11_n_869 = (mul_72_11_n_475 ^ (mul_72_11_n_434 ^ mul_72_11_n_752));
 assign mul_72_11_n_866 = ((mul_72_11_n_755 & mul_72_11_n_405) | ((mul_72_11_n_405 & mul_72_11_n_479)
    | (mul_72_11_n_479 & mul_72_11_n_755)));
 assign mul_72_11_n_867 = (mul_72_11_n_405 ^ (mul_72_11_n_479 ^ mul_72_11_n_755));
 assign mul_72_11_n_864 = ((mul_72_11_n_740 & mul_72_11_n_474) | ((mul_72_11_n_474 & mul_72_11_n_453)
    | (mul_72_11_n_453 & mul_72_11_n_740)));
 assign mul_72_11_n_865 = (mul_72_11_n_474 ^ (mul_72_11_n_453 ^ mul_72_11_n_740));
 assign mul_72_11_n_862 = ((mul_72_11_n_760 & mul_72_11_n_490) | ((mul_72_11_n_490 & mul_72_11_n_467)
    | (mul_72_11_n_467 & mul_72_11_n_760)));
 assign mul_72_11_n_863 = (mul_72_11_n_490 ^ (mul_72_11_n_467 ^ mul_72_11_n_760));
 assign mul_72_11_n_861 = ~(mul_72_11_n_852 & ~mul_72_11_n_851);
 assign mul_72_11_n_860 = ~(mul_72_11_n_836 & mul_72_11_n_767);
 assign mul_72_11_n_874 = ~(mul_72_11_n_851 | mul_72_11_n_836);
 assign mul_72_11_n_858 = ~mul_72_11_n_857;
 assign {out1[4]} = ~(mul_72_11_n_794 ^ mul_72_11_n_832);
 assign mul_72_11_n_855 = ~(mul_72_11_n_693 ^ mul_72_11_n_803);
 assign mul_72_11_n_859 = ~(mul_72_11_n_854 | mul_72_11_n_833);
 assign mul_72_11_n_857 = (mul_72_11_n_854 & mul_72_11_n_833);
 assign mul_72_11_n_849 = ((mul_72_11_n_781 & mul_72_11_n_599) | ((mul_72_11_n_599 & mul_72_11_n_723)
    | (mul_72_11_n_723 & mul_72_11_n_781)));
 assign mul_72_11_n_850 = (mul_72_11_n_599 ^ (mul_72_11_n_723 ^ mul_72_11_n_781));
 assign mul_72_11_n_847 = ((mul_72_11_n_753 & mul_72_11_n_594) | ((mul_72_11_n_594 & mul_72_11_n_721)
    | (mul_72_11_n_721 & mul_72_11_n_753)));
 assign mul_72_11_n_848 = (mul_72_11_n_594 ^ (mul_72_11_n_721 ^ mul_72_11_n_753));
 assign mul_72_11_n_845 = ((mul_72_11_n_777 & mul_72_11_n_380) | ((mul_72_11_n_380 & mul_72_11_n_430)
    | (mul_72_11_n_430 & mul_72_11_n_777)));
 assign mul_72_11_n_846 = (mul_72_11_n_380 ^ (mul_72_11_n_430 ^ mul_72_11_n_777));
 assign mul_72_11_n_843 = ((mul_72_11_n_779 & mul_72_11_n_381) | ((mul_72_11_n_381 & mul_72_11_n_425)
    | (mul_72_11_n_425 & mul_72_11_n_779)));
 assign mul_72_11_n_844 = (mul_72_11_n_381 ^ (mul_72_11_n_425 ^ mul_72_11_n_779));
 assign mul_72_11_n_853 = ((mul_72_11_n_787 & mul_72_11_n_406) | ((mul_72_11_n_406 & mul_72_11_n_423)
    | (mul_72_11_n_423 & mul_72_11_n_787)));
 assign mul_72_11_n_854 = (mul_72_11_n_406 ^ (mul_72_11_n_423 ^ mul_72_11_n_787));
 assign mul_72_11_n_841 = ((mul_72_11_n_785 & mul_72_11_n_593) | ((mul_72_11_n_593 & mul_72_11_n_431)
    | (mul_72_11_n_431 & mul_72_11_n_785)));
 assign mul_72_11_n_842 = (mul_72_11_n_593 ^ (mul_72_11_n_431 ^ mul_72_11_n_785));
 assign mul_72_11_n_839 = ((mul_72_11_n_775 & mul_72_11_n_555) | ((mul_72_11_n_555 & mul_72_11_n_704)
    | (mul_72_11_n_704 & mul_72_11_n_775)));
 assign mul_72_11_n_840 = (mul_72_11_n_555 ^ (mul_72_11_n_704 ^ mul_72_11_n_775));
 assign mul_72_11_n_837 = ((mul_72_11_n_761 & mul_72_11_n_563) | ((mul_72_11_n_563 & mul_72_11_n_698)
    | (mul_72_11_n_698 & mul_72_11_n_761)));
 assign mul_72_11_n_838 = (mul_72_11_n_563 ^ (mul_72_11_n_698 ^ mul_72_11_n_761));
 assign mul_72_11_n_852 = ~(mul_72_11_n_834 & mul_72_11_n_764);
 assign mul_72_11_n_851 = ~(mul_72_11_n_834 | mul_72_11_n_764);
 assign mul_72_11_n_836 = ~(mul_72_11_n_832 & ~mul_72_11_n_792);
 assign mul_72_11_n_835 = ~(mul_72_11_n_793 ^ mul_72_11_n_487);
 assign mul_72_11_n_830 = ((mul_72_11_n_705 & mul_72_11_n_602) | ((mul_72_11_n_602 & mul_72_11_n_439)
    | (mul_72_11_n_439 & mul_72_11_n_705)));
 assign mul_72_11_n_831 = (mul_72_11_n_602 ^ (mul_72_11_n_439 ^ mul_72_11_n_705));
 assign mul_72_11_n_828 = ((mul_72_11_n_708 & mul_72_11_n_462) | ((mul_72_11_n_462 & mul_72_11_n_601)
    | (mul_72_11_n_601 & mul_72_11_n_708)));
 assign mul_72_11_n_829 = (mul_72_11_n_462 ^ (mul_72_11_n_601 ^ mul_72_11_n_708));
 assign mul_72_11_n_826 = ((mul_72_11_n_719 & mul_72_11_n_459) | ((mul_72_11_n_459 & mul_72_11_n_600)
    | (mul_72_11_n_600 & mul_72_11_n_719)));
 assign mul_72_11_n_827 = (mul_72_11_n_459 ^ (mul_72_11_n_600 ^ mul_72_11_n_719));
 assign mul_72_11_n_824 = ((mul_72_11_n_701 & mul_72_11_n_556) | ((mul_72_11_n_556 & mul_72_11_n_441)
    | (mul_72_11_n_441 & mul_72_11_n_701)));
 assign mul_72_11_n_825 = (mul_72_11_n_556 ^ (mul_72_11_n_441 ^ mul_72_11_n_701));
 assign mul_72_11_n_822 = ((mul_72_11_n_707 & mul_72_11_n_597) | ((mul_72_11_n_597 & mul_72_11_n_446)
    | (mul_72_11_n_446 & mul_72_11_n_707)));
 assign mul_72_11_n_823 = (mul_72_11_n_597 ^ (mul_72_11_n_446 ^ mul_72_11_n_707));
 assign mul_72_11_n_820 = ((mul_72_11_n_703 & mul_72_11_n_592) | ((mul_72_11_n_592 & mul_72_11_n_422)
    | (mul_72_11_n_422 & mul_72_11_n_703)));
 assign mul_72_11_n_821 = (mul_72_11_n_592 ^ (mul_72_11_n_422 ^ mul_72_11_n_703));
 assign mul_72_11_n_818 = ((mul_72_11_n_713 & mul_72_11_n_458) | ((mul_72_11_n_458 & mul_72_11_n_596)
    | (mul_72_11_n_596 & mul_72_11_n_713)));
 assign mul_72_11_n_819 = (mul_72_11_n_458 ^ (mul_72_11_n_596 ^ mul_72_11_n_713));
 assign mul_72_11_n_816 = ((mul_72_11_n_720 & mul_72_11_n_598) | ((mul_72_11_n_598 & mul_72_11_n_436)
    | (mul_72_11_n_436 & mul_72_11_n_720)));
 assign mul_72_11_n_817 = (mul_72_11_n_598 ^ (mul_72_11_n_436 ^ mul_72_11_n_720));
 assign mul_72_11_n_814 = ((mul_72_11_n_714 & mul_72_11_n_588) | ((mul_72_11_n_588 & mul_72_11_n_432)
    | (mul_72_11_n_432 & mul_72_11_n_714)));
 assign mul_72_11_n_815 = (mul_72_11_n_588 ^ (mul_72_11_n_432 ^ mul_72_11_n_714));
 assign mul_72_11_n_812 = ((mul_72_11_n_722 & mul_72_11_n_561) | ((mul_72_11_n_561 & mul_72_11_n_427)
    | (mul_72_11_n_427 & mul_72_11_n_722)));
 assign mul_72_11_n_813 = (mul_72_11_n_561 ^ (mul_72_11_n_427 ^ mul_72_11_n_722));
 assign mul_72_11_n_810 = ((mul_72_11_n_716 & mul_72_11_n_670) | ((mul_72_11_n_670 & mul_72_11_n_424)
    | (mul_72_11_n_424 & mul_72_11_n_716)));
 assign mul_72_11_n_811 = (mul_72_11_n_670 ^ (mul_72_11_n_424 ^ mul_72_11_n_716));
 assign mul_72_11_n_833 = ((mul_72_11_n_712 & mul_72_11_n_444) | ((mul_72_11_n_444 & mul_72_11_n_573)
    | (mul_72_11_n_573 & mul_72_11_n_712)));
 assign mul_72_11_n_834 = (mul_72_11_n_444 ^ (mul_72_11_n_573 ^ mul_72_11_n_712));
 assign mul_72_11_n_832 = ((mul_72_11_n_746 & mul_72_11_n_621) | ((mul_72_11_n_621 & mul_72_11_n_710)
    | (mul_72_11_n_710 & mul_72_11_n_746)));
 assign {out1[3]} = (mul_72_11_n_621 ^ (mul_72_11_n_710 ^ mul_72_11_n_746));
 assign mul_72_11_n_807 = ((mul_72_11_n_718 & mul_72_11_n_402) | ((mul_72_11_n_402 & mul_72_11_n_426)
    | (mul_72_11_n_426 & mul_72_11_n_718)));
 assign mul_72_11_n_808 = (mul_72_11_n_402 ^ (mul_72_11_n_426 ^ mul_72_11_n_718));
 assign mul_72_11_n_805 = ((mul_72_11_n_709 & mul_72_11_n_560) | ((mul_72_11_n_560 & mul_72_11_n_437)
    | (mul_72_11_n_437 & mul_72_11_n_709)));
 assign mul_72_11_n_806 = (mul_72_11_n_560 ^ (mul_72_11_n_437 ^ mul_72_11_n_709));
 assign mul_72_11_n_803 = ((mul_72_11_n_702 & mul_72_11_n_466) | ((mul_72_11_n_466 & mul_72_11_n_566)
    | (mul_72_11_n_566 & mul_72_11_n_702)));
 assign mul_72_11_n_804 = (mul_72_11_n_466 ^ (mul_72_11_n_566 ^ mul_72_11_n_702));
 assign mul_72_11_n_801 = ((mul_72_11_n_699 & mul_72_11_n_562) | ((mul_72_11_n_562 & mul_72_11_n_442)
    | (mul_72_11_n_442 & mul_72_11_n_699)));
 assign mul_72_11_n_802 = (mul_72_11_n_562 ^ (mul_72_11_n_442 ^ mul_72_11_n_699));
 assign mul_72_11_n_799 = ((mul_72_11_n_706 & mul_72_11_n_469) | ((mul_72_11_n_469 & mul_72_11_n_587)
    | (mul_72_11_n_587 & mul_72_11_n_706)));
 assign mul_72_11_n_800 = (mul_72_11_n_469 ^ (mul_72_11_n_587 ^ mul_72_11_n_706));
 assign mul_72_11_n_797 = ((mul_72_11_n_724 & mul_72_11_n_595) | ((mul_72_11_n_595 & mul_72_11_n_433)
    | (mul_72_11_n_433 & mul_72_11_n_724)));
 assign mul_72_11_n_798 = (mul_72_11_n_595 ^ (mul_72_11_n_433 ^ mul_72_11_n_724));
 assign mul_72_11_n_795 = ((mul_72_11_n_728 & mul_72_11_n_500) | ((mul_72_11_n_500 & mul_72_11_n_659)
    | (mul_72_11_n_659 & mul_72_11_n_728)));
 assign mul_72_11_n_796 = (mul_72_11_n_500 ^ (mul_72_11_n_659 ^ mul_72_11_n_728));
 assign mul_72_11_n_794 = ~(mul_72_11_n_767 & ~mul_72_11_n_792);
 assign mul_72_11_n_793 = ~(mul_72_11_n_488 ^ mul_72_11_n_738);
 assign mul_72_11_n_790 = ((mul_72_11_n_680 & mul_72_11_n_496) | ((mul_72_11_n_496 & mul_72_11_n_645)
    | (mul_72_11_n_645 & mul_72_11_n_680)));
 assign mul_72_11_n_791 = (mul_72_11_n_496 ^ (mul_72_11_n_645 ^ mul_72_11_n_680));
 assign mul_72_11_n_788 = ((mul_72_11_n_675 & mul_72_11_n_384) | ((mul_72_11_n_384 & mul_72_11_n_571)
    | (mul_72_11_n_571 & mul_72_11_n_675)));
 assign mul_72_11_n_789 = (mul_72_11_n_384 ^ (mul_72_11_n_571 ^ mul_72_11_n_675));
 assign mul_72_11_n_786 = ((mul_72_11_n_711 & mul_72_11_n_523) | ((mul_72_11_n_523 & mul_72_11_n_584)
    | (mul_72_11_n_584 & mul_72_11_n_711)));
 assign mul_72_11_n_787 = (mul_72_11_n_523 ^ (mul_72_11_n_584 ^ mul_72_11_n_711));
 assign mul_72_11_n_784 = ((mul_72_11_n_717 & mul_72_11_n_499) | ((mul_72_11_n_499 & mul_72_11_n_568)
    | (mul_72_11_n_568 & mul_72_11_n_717)));
 assign mul_72_11_n_785 = (mul_72_11_n_499 ^ (mul_72_11_n_568 ^ mul_72_11_n_717));
 assign mul_72_11_n_782 = ((mul_72_11_n_483 & mul_72_11_n_525) | ((mul_72_11_n_525 & mul_72_11_n_572)
    | (mul_72_11_n_572 & mul_72_11_n_483)));
 assign mul_72_11_n_783 = (mul_72_11_n_525 ^ (mul_72_11_n_572 ^ mul_72_11_n_483));
 assign mul_72_11_n_780 = ((mul_72_11_n_485 & mul_72_11_n_501) | ((mul_72_11_n_501 & mul_72_11_n_580)
    | (mul_72_11_n_580 & mul_72_11_n_485)));
 assign mul_72_11_n_781 = (mul_72_11_n_501 ^ (mul_72_11_n_580 ^ mul_72_11_n_485));
 assign mul_72_11_n_778 = ((mul_72_11_n_700 & mul_72_11_n_518) | ((mul_72_11_n_518 & mul_72_11_n_564)
    | (mul_72_11_n_564 & mul_72_11_n_700)));
 assign mul_72_11_n_779 = (mul_72_11_n_518 ^ (mul_72_11_n_564 ^ mul_72_11_n_700));
 assign mul_72_11_n_776 = ((mul_72_11_n_715 & mul_72_11_n_521) | ((mul_72_11_n_521 & mul_72_11_n_565)
    | (mul_72_11_n_565 & mul_72_11_n_715)));
 assign mul_72_11_n_777 = (mul_72_11_n_521 ^ (mul_72_11_n_565 ^ mul_72_11_n_715));
 assign mul_72_11_n_774 = ((mul_72_11_n_484 & mul_72_11_n_489) | ((mul_72_11_n_489 & mul_72_11_n_579)
    | (mul_72_11_n_579 & mul_72_11_n_484)));
 assign mul_72_11_n_775 = (mul_72_11_n_489 ^ (mul_72_11_n_579 ^ mul_72_11_n_484));
 assign mul_72_11_n_772 = ((mul_72_11_n_530 & mul_72_11_n_656) | ((mul_72_11_n_656 & mul_72_11_n_642)
    | (mul_72_11_n_642 & mul_72_11_n_530)));
 assign mul_72_11_n_773 = (mul_72_11_n_656 ^ (mul_72_11_n_642 ^ mul_72_11_n_530));
 assign mul_72_11_n_770 = ((mul_72_11_n_674 & mul_72_11_n_409) | ((mul_72_11_n_409 & mul_72_11_n_627)
    | (mul_72_11_n_627 & mul_72_11_n_674)));
 assign mul_72_11_n_771 = (mul_72_11_n_409 ^ (mul_72_11_n_627 ^ mul_72_11_n_674));
 assign mul_72_11_n_768 = ((mul_72_11_n_682 & mul_72_11_n_508) | ((mul_72_11_n_508 & mul_72_11_n_651)
    | (mul_72_11_n_651 & mul_72_11_n_682)));
 assign mul_72_11_n_769 = (mul_72_11_n_508 ^ (mul_72_11_n_651 ^ mul_72_11_n_682));
 assign mul_72_11_n_792 = ~(mul_72_11_n_765 | mul_72_11_n_725);
 assign mul_72_11_n_766 = ~(mul_72_11_n_685 ^ mul_72_11_n_726);
 assign mul_72_11_n_767 = ~(mul_72_11_n_765 & mul_72_11_n_725);
 assign mul_72_11_n_762 = ((mul_72_11_n_620 & mul_72_11_n_385) | ((mul_72_11_n_385 & mul_72_11_n_630)
    | (mul_72_11_n_630 & mul_72_11_n_620)));
 assign mul_72_11_n_763 = (mul_72_11_n_385 ^ (mul_72_11_n_630 ^ mul_72_11_n_620));
 assign mul_72_11_n_760 = ((mul_72_11_n_537 & mul_72_11_n_445) | ((mul_72_11_n_445 & mul_72_11_n_582)
    | (mul_72_11_n_582 & mul_72_11_n_537)));
 assign mul_72_11_n_761 = (mul_72_11_n_445 ^ (mul_72_11_n_582 ^ mul_72_11_n_537));
 assign mul_72_11_n_758 = ((mul_72_11_n_603 & mul_72_11_n_401) | ((mul_72_11_n_401 & mul_72_11_n_636)
    | (mul_72_11_n_636 & mul_72_11_n_603)));
 assign mul_72_11_n_759 = (mul_72_11_n_401 ^ (mul_72_11_n_636 ^ mul_72_11_n_603));
 assign mul_72_11_n_756 = ((mul_72_11_n_677 & mul_72_11_n_505) | ((mul_72_11_n_505 & mul_72_11_n_494)
    | (mul_72_11_n_494 & mul_72_11_n_677)));
 assign mul_72_11_n_757 = (mul_72_11_n_505 ^ (mul_72_11_n_494 ^ mul_72_11_n_677));
 assign mul_72_11_n_754 = ((mul_72_11_n_616 & mul_72_11_n_438) | ((mul_72_11_n_438 & mul_72_11_n_504)
    | (mul_72_11_n_504 & mul_72_11_n_616)));
 assign mul_72_11_n_755 = (mul_72_11_n_438 ^ (mul_72_11_n_504 ^ mul_72_11_n_616));
 assign mul_72_11_n_764 = ((mul_72_11_n_615 & mul_72_11_n_383) | ((mul_72_11_n_383 & mul_72_11_n_520)
    | (mul_72_11_n_520 & mul_72_11_n_615)));
 assign mul_72_11_n_765 = (mul_72_11_n_383 ^ (mul_72_11_n_520 ^ mul_72_11_n_615));
 assign mul_72_11_n_752 = ((mul_72_11_n_611 & mul_72_11_n_428) | ((mul_72_11_n_428 & mul_72_11_n_510)
    | (mul_72_11_n_510 & mul_72_11_n_611)));
 assign mul_72_11_n_753 = (mul_72_11_n_428 ^ (mul_72_11_n_510 ^ mul_72_11_n_611));
 assign mul_72_11_n_750 = ((mul_72_11_n_546 & mul_72_11_n_658) | ((mul_72_11_n_658 & mul_72_11_n_626)
    | (mul_72_11_n_626 & mul_72_11_n_546)));
 assign mul_72_11_n_751 = (mul_72_11_n_658 ^ (mul_72_11_n_626 ^ mul_72_11_n_546));
 assign mul_72_11_n_748 = ((mul_72_11_n_527 & mul_72_11_n_583) | ((mul_72_11_n_583 & mul_72_11_n_443)
    | (mul_72_11_n_443 & mul_72_11_n_527)));
 assign mul_72_11_n_749 = (mul_72_11_n_583 ^ (mul_72_11_n_443 ^ mul_72_11_n_527));
 assign mul_72_11_n_746 = ((mul_72_11_n_689 & mul_72_11_n_407) | ((mul_72_11_n_407 & mul_72_11_n_552)
    | (mul_72_11_n_552 & mul_72_11_n_689)));
 assign {out1[2]} = (mul_72_11_n_407 ^ (mul_72_11_n_552 ^ mul_72_11_n_689));
 assign mul_72_11_n_744 = ((mul_72_11_n_679 & mul_72_11_n_509) | ((mul_72_11_n_509 & mul_72_11_n_498)
    | (mul_72_11_n_498 & mul_72_11_n_679)));
 assign mul_72_11_n_745 = (mul_72_11_n_509 ^ (mul_72_11_n_498 ^ mul_72_11_n_679));
 assign mul_72_11_n_742 = ((mul_72_11_n_542 & mul_72_11_n_515) | ((mul_72_11_n_515 & mul_72_11_n_493)
    | (mul_72_11_n_493 & mul_72_11_n_542)));
 assign mul_72_11_n_743 = (mul_72_11_n_515 ^ (mul_72_11_n_493 ^ mul_72_11_n_542));
 assign mul_72_11_n_740 = ((mul_72_11_n_676 & mul_72_11_n_429) | ((mul_72_11_n_429 & mul_72_11_n_524)
    | (mul_72_11_n_524 & mul_72_11_n_676)));
 assign mul_72_11_n_741 = (mul_72_11_n_429 ^ (mul_72_11_n_524 ^ mul_72_11_n_676));
 assign mul_72_11_n_738 = ((mul_72_11_n_544 & mul_72_11_n_526) | ((mul_72_11_n_526 & mul_72_11_n_664)
    | (mul_72_11_n_664 & mul_72_11_n_544)));
 assign mul_72_11_n_739 = (mul_72_11_n_526 ^ (mul_72_11_n_664 ^ mul_72_11_n_544));
 assign mul_72_11_n_736 = ((mul_72_11_n_605 & mul_72_11_n_649) | ((mul_72_11_n_649 & mul_72_11_n_634)
    | (mul_72_11_n_634 & mul_72_11_n_605)));
 assign mul_72_11_n_737 = (mul_72_11_n_649 ^ (mul_72_11_n_634 ^ mul_72_11_n_605));
 assign mul_72_11_n_734 = ((mul_72_11_n_681 & mul_72_11_n_648) | ((mul_72_11_n_648 & mul_72_11_n_517)
    | (mul_72_11_n_517 & mul_72_11_n_681)));
 assign mul_72_11_n_735 = (mul_72_11_n_648 ^ (mul_72_11_n_517 ^ mul_72_11_n_681));
 assign mul_72_11_n_732 = ((mul_72_11_n_486 & mul_72_11_n_404) | ((mul_72_11_n_404 & mul_72_11_n_471)
    | (mul_72_11_n_471 & mul_72_11_n_486)));
 assign mul_72_11_n_733 = (mul_72_11_n_404 ^ (mul_72_11_n_471 ^ mul_72_11_n_486));
 assign mul_72_11_n_730 = ((mul_72_11_n_538 & mul_72_11_n_666) | ((mul_72_11_n_666 & mul_72_11_n_513)
    | (mul_72_11_n_513 & mul_72_11_n_538)));
 assign mul_72_11_n_731 = (mul_72_11_n_666 ^ (mul_72_11_n_513 ^ mul_72_11_n_538));
 assign mul_72_11_n_728 = ((mul_72_11_n_482 & mul_72_11_n_379) | ((mul_72_11_n_379 & mul_72_11_n_450)
    | (mul_72_11_n_450 & mul_72_11_n_482)));
 assign mul_72_11_n_729 = (mul_72_11_n_379 ^ (mul_72_11_n_450 ^ mul_72_11_n_482));
 assign mul_72_11_n_727 = ~(mul_72_11_n_692 ^ mul_72_11_n_553);
 assign mul_72_11_n_726 = ~(mul_72_11_n_696 ^ mul_72_11_n_695);
 assign mul_72_11_n_723 = (mul_72_11_n_613 & mul_72_11_n_532);
 assign mul_72_11_n_724 = (mul_72_11_n_613 ^ mul_72_11_n_532);
 assign mul_72_11_n_721 = (mul_72_11_n_606 & mul_72_11_n_533);
 assign mul_72_11_n_722 = (mul_72_11_n_606 ^ mul_72_11_n_533);
 assign mul_72_11_n_719 = (mul_72_11_n_614 & mul_72_11_n_545);
 assign mul_72_11_n_720 = (mul_72_11_n_614 ^ mul_72_11_n_545);
 assign mul_72_11_n_717 = (mul_72_11_n_609 & mul_72_11_n_540);
 assign mul_72_11_n_718 = (mul_72_11_n_609 ^ mul_72_11_n_540);
 assign mul_72_11_n_715 = (mul_72_11_n_607 & mul_72_11_n_539);
 assign mul_72_11_n_716 = (mul_72_11_n_607 ^ mul_72_11_n_539);
 assign mul_72_11_n_713 = (mul_72_11_n_612 & mul_72_11_n_535);
 assign mul_72_11_n_714 = (mul_72_11_n_612 ^ mul_72_11_n_535);
 assign mul_72_11_n_711 = (mul_72_11_n_529 & mul_72_11_n_619);
 assign mul_72_11_n_712 = (mul_72_11_n_529 ^ mul_72_11_n_619);
 assign mul_72_11_n_725 = (mul_72_11_n_531 & mul_72_11_n_678);
 assign mul_72_11_n_710 = (mul_72_11_n_531 ^ mul_72_11_n_678);
 assign mul_72_11_n_708 = (mul_72_11_n_608 & mul_72_11_n_543);
 assign mul_72_11_n_709 = (mul_72_11_n_608 ^ mul_72_11_n_543);
 assign mul_72_11_n_706 = (mul_72_11_n_610 & mul_72_11_n_534);
 assign mul_72_11_n_707 = (mul_72_11_n_610 ^ mul_72_11_n_534);
 assign mul_72_11_n_704 = (mul_72_11_n_617 & mul_72_11_n_547);
 assign mul_72_11_n_705 = (mul_72_11_n_617 ^ mul_72_11_n_547);
 assign mul_72_11_n_702 = (mul_72_11_n_673 & mul_72_11_n_528);
 assign mul_72_11_n_703 = (mul_72_11_n_673 ^ mul_72_11_n_528);
 assign mul_72_11_n_700 = (mul_72_11_n_604 & mul_72_11_n_536);
 assign mul_72_11_n_701 = (mul_72_11_n_604 ^ mul_72_11_n_536);
 assign mul_72_11_n_698 = (mul_72_11_n_618 & mul_72_11_n_541);
 assign mul_72_11_n_699 = (mul_72_11_n_618 ^ mul_72_11_n_541);
 assign mul_72_11_n_697 = ~(mul_72_11_n_690 ^ mul_72_11_n_688);
 assign mul_72_11_n_696 = ~(mul_72_11_n_622 ^ mul_72_11_n_551);
 assign mul_72_11_n_695 = ~(mul_72_11_n_548 ^ mul_72_11_n_686);
 assign mul_72_11_n_694 = ~(mul_72_11_n_12 ^ mul_72_11_n_15);
 assign mul_72_11_n_693 = ~(mul_72_11_n_687 ^ mul_72_11_n_14);
 assign mul_72_11_n_692 = ~(mul_72_11_n_683 ^ mul_72_11_n_684);
 assign {out1[1]} = ~(mul_72_11_n_689 | (mul_72_11_n_554 & mul_72_11_n_330));
 assign mul_72_11_n_690 = ~(mul_72_11_n_549 ^ mul_72_11_n_550);
 assign mul_72_11_n_688 = ~((mul_72_11_n_421 & mul_72_11_n_275) | (mul_72_11_n_395 & mul_72_11_n_248));
 assign mul_72_11_n_687 = ~(mul_72_11_n_408 & (n_397 & (mul_72_11_n_55 | mul_72_11_n_37)));
 assign mul_72_11_n_686 = ~((mul_72_11_n_13 | mul_72_11_n_364) & (mul_72_11_n_249 | mul_72_11_n_247));
 assign mul_72_11_n_685 = ~((mul_72_11_n_413 & mul_72_11_n_295) | (mul_72_11_n_256 & mul_72_11_n_222));
 assign mul_72_11_n_684 = ~((mul_72_11_n_419 & mul_72_11_n_177) | (mul_72_11_n_396 & mul_72_11_n_79));
 assign mul_72_11_n_683 = ~((mul_72_11_n_417 & mul_72_11_n_106) | (mul_72_11_n_397 & mul_72_11_n_71));
 assign mul_72_11_n_682 = ~((mul_72_11_n_416 | mul_72_11_n_99) & (mul_72_11_n_261 | mul_72_11_n_90));
 assign mul_72_11_n_681 = ~((mul_72_11_n_416 | mul_72_11_n_90) & (mul_72_11_n_261 | mul_72_11_n_91));
 assign mul_72_11_n_680 = ~((mul_72_11_n_416 | mul_72_11_n_73) & (mul_72_11_n_261 | mul_72_11_n_109));
 assign mul_72_11_n_679 = ~((mul_72_11_n_415 | mul_72_11_n_193) & (mul_72_11_n_257 | mul_72_11_n_194));
 assign mul_72_11_n_677 = ~((mul_72_11_n_415 | mul_72_11_n_160) & (mul_72_11_n_257 | mul_72_11_n_161));
 assign mul_72_11_n_676 = ~((mul_72_11_n_13 | mul_72_11_n_371) & (mul_72_11_n_249 | mul_72_11_n_335));
 assign mul_72_11_n_675 = ~((mul_72_11_n_414 | mul_72_11_n_125) & (mul_72_11_n_399 | mul_72_11_n_136));
 assign mul_72_11_n_674 = ~((mul_72_11_n_414 | mul_72_11_n_146) & (mul_72_11_n_399 | mul_72_11_n_271));
 assign mul_72_11_n_673 = ~((mul_72_11_n_13 | mul_72_11_n_335) & (mul_72_11_n_249 | mul_72_11_n_359));
 assign mul_72_11_n_668 = ~((mul_72_11_n_420 | mul_72_11_n_225) & (mul_72_11_n_264 | mul_72_11_n_282));
 assign mul_72_11_n_667 = ~((mul_72_11_n_416 | mul_72_11_n_92) & (mul_72_11_n_261 | mul_72_11_n_105));
 assign mul_72_11_n_666 = ~((mul_72_11_n_416 | mul_72_11_n_93) & (mul_72_11_n_261 | mul_72_11_n_92));
 assign mul_72_11_n_664 = ~((mul_72_11_n_13 | mul_72_11_n_359) & (mul_72_11_n_249 | mul_72_11_n_364));
 assign mul_72_11_n_663 = ~((mul_72_11_n_420 | mul_72_11_n_282) & (mul_72_11_n_264 | mul_72_11_n_274));
 assign mul_72_11_n_662 = ~((mul_72_11_n_416 | mul_72_11_n_91) & (mul_72_11_n_261 | mul_72_11_n_93));
 assign mul_72_11_n_661 = ~((mul_72_11_n_416 | mul_72_11_n_98) & (mul_72_11_n_261 | mul_72_11_n_99));
 assign mul_72_11_n_660 = ~((mul_72_11_n_416 | mul_72_11_n_109) & (mul_72_11_n_261 | mul_72_11_n_98));
 assign mul_72_11_n_659 = ~((mul_72_11_n_415 | mul_72_11_n_126) & (mul_72_11_n_257 | mul_72_11_n_127));
 assign mul_72_11_n_658 = ~((mul_72_11_n_415 | mul_72_11_n_127) & (mul_72_11_n_257 | mul_72_11_n_140));
 assign mul_72_11_n_657 = ~((mul_72_11_n_415 | mul_72_11_n_84) & (mul_72_11_n_257 | mul_72_11_n_367));
 assign mul_72_11_n_656 = ~((mul_72_11_n_415 | mul_72_11_n_116) & (mul_72_11_n_257 | mul_72_11_n_126));
 assign mul_72_11_n_689 = ~(mul_72_11_n_554 | mul_72_11_n_330);
 assign mul_72_11_n_655 = ~((mul_72_11_n_415 | mul_72_11_n_194) & (mul_72_11_n_257 | mul_72_11_n_85));
 assign mul_72_11_n_652 = ~((mul_72_11_n_415 | mul_72_11_n_115) & (mul_72_11_n_257 | mul_72_11_n_116));
 assign mul_72_11_n_651 = ~((mul_72_11_n_415 | mul_72_11_n_161) & (mul_72_11_n_257 | mul_72_11_n_193));
 assign mul_72_11_n_650 = ~((mul_72_11_n_415 | mul_72_11_n_103) & (mul_72_11_n_257 | mul_72_11_n_115));
 assign mul_72_11_n_649 = ~((mul_72_11_n_415 | mul_72_11_n_75) & (mul_72_11_n_257 | mul_72_11_n_103));
 assign mul_72_11_n_648 = ~((mul_72_11_n_418 | mul_72_11_n_221) & (mul_72_11_n_263 | mul_72_11_n_205));
 assign mul_72_11_n_647 = ~((mul_72_11_n_415 | mul_72_11_n_85) & (mul_72_11_n_257 | mul_72_11_n_84));
 assign mul_72_11_n_646 = ~((mul_72_11_n_415 | mul_72_11_n_141) & (mul_72_11_n_257 | mul_72_11_n_160));
 assign mul_72_11_n_645 = ~((mul_72_11_n_415 | mul_72_11_n_140) & (mul_72_11_n_257 | mul_72_11_n_141));
 assign mul_72_11_n_644 = ~((mul_72_11_n_414 | mul_72_11_n_271) & (mul_72_11_n_399 | mul_72_11_n_272));
 assign mul_72_11_n_643 = ~((mul_72_11_n_414 | mul_72_11_n_155) & (mul_72_11_n_399 | mul_72_11_n_181));
 assign mul_72_11_n_642 = ~((mul_72_11_n_414 | mul_72_11_n_137) & (mul_72_11_n_399 | mul_72_11_n_156));
 assign mul_72_11_n_641 = ~((mul_72_11_n_414 | mul_72_11_n_156) & (mul_72_11_n_399 | mul_72_11_n_155));
 assign mul_72_11_n_640 = ~((mul_72_11_n_414 | mul_72_11_n_148) & (mul_72_11_n_399 | mul_72_11_n_146));
 assign mul_72_11_n_639 = ~((mul_72_11_n_414 | mul_72_11_n_136) & (mul_72_11_n_399 | mul_72_11_n_137));
 assign mul_72_11_n_638 = ~((mul_72_11_n_418 | mul_72_11_n_205) & (mul_72_11_n_263 | mul_72_11_n_190));
 assign mul_72_11_n_637 = ~((mul_72_11_n_418 | mul_72_11_n_190) & (mul_72_11_n_263 | mul_72_11_n_189));
 assign mul_72_11_n_636 = ~((mul_72_11_n_414 | mul_72_11_n_210) & (mul_72_11_n_399 | mul_72_11_n_148));
 assign mul_72_11_n_635 = ~((mul_72_11_n_418 | mul_72_11_n_189) & (mul_72_11_n_263 | mul_72_11_n_176));
 assign mul_72_11_n_634 = ~((mul_72_11_n_414 | mul_72_11_n_124) & (mul_72_11_n_399 | mul_72_11_n_125));
 assign mul_72_11_n_633 = ~((mul_72_11_n_414 | mul_72_11_n_211) & (mul_72_11_n_399 | mul_72_11_n_210));
 assign mul_72_11_n_632 = ~((mul_72_11_n_414 | mul_72_11_n_117) & (mul_72_11_n_399 | mul_72_11_n_124));
 assign mul_72_11_n_631 = ~((mul_72_11_n_414 | mul_72_11_n_74) & (mul_72_11_n_399 | mul_72_11_n_117));
 assign mul_72_11_n_630 = ~((mul_72_11_n_414 | mul_72_11_n_272) & (mul_72_11_n_399 | mul_72_11_n_296));
 assign mul_72_11_n_629 = ~((mul_72_11_n_414 | mul_72_11_n_181) & (mul_72_11_n_399 | mul_72_11_n_182));
 assign mul_72_11_n_628 = ~((mul_72_11_n_414 | mul_72_11_n_182) & (mul_72_11_n_399 | mul_72_11_n_211));
 assign mul_72_11_n_627 = ~((mul_72_11_n_412 | mul_72_11_n_279) & (mul_72_11_n_255 | mul_72_11_n_303));
 assign mul_72_11_n_626 = ~((mul_72_11_n_412 | mul_72_11_n_197) & (mul_72_11_n_255 | mul_72_11_n_219));
 assign mul_72_11_n_625 = ~((mul_72_11_n_412 | mul_72_11_n_121) & (mul_72_11_n_255 | mul_72_11_n_134));
 assign mul_72_11_n_624 = ~((mul_72_11_n_412 | mul_72_11_n_198) & (mul_72_11_n_255 | mul_72_11_n_197));
 assign mul_72_11_n_623 = ~((mul_72_11_n_412 | mul_72_11_n_172) & (mul_72_11_n_255 | mul_72_11_n_198));
 assign mul_72_11_n_622 = ~((mul_72_11_n_410 & mul_72_11_n_365) | (mul_72_11_n_394 & mul_72_11_n_231));
 assign mul_72_11_n_621 = ~((mul_72_11_n_13 | mul_72_11_n_66) & (mul_72_11_n_249 | mul_72_11_n_162));
 assign mul_72_11_n_620 = ~((mul_72_11_n_412 | mul_72_11_n_302) & (mul_72_11_n_255 | mul_72_11_n_320));
 assign mul_72_11_n_618 = ~((mul_72_11_n_13 | mul_72_11_n_315) & (mul_72_11_n_249 | mul_72_11_n_316));
 assign mul_72_11_n_617 = ~((mul_72_11_n_13 | mul_72_11_n_301) & (mul_72_11_n_249 | mul_72_11_n_300));
 assign mul_72_11_n_616 = ~((mul_72_11_n_13 | mul_72_11_n_283) & (mul_72_11_n_249 | mul_72_11_n_301));
 assign mul_72_11_n_615 = ~((mul_72_11_n_13 | mul_72_11_n_162) & (mul_72_11_n_249 | mul_72_11_n_180));
 assign mul_72_11_n_614 = ~((mul_72_11_n_13 | mul_72_11_n_284) & (mul_72_11_n_249 | mul_72_11_n_283));
 assign mul_72_11_n_613 = ~((mul_72_11_n_13 | mul_72_11_n_343) & (mul_72_11_n_249 | mul_72_11_n_344));
 assign mul_72_11_n_612 = ~((mul_72_11_n_13 | mul_72_11_n_360) & (mul_72_11_n_249 | mul_72_11_n_291));
 assign mul_72_11_n_611 = ~((mul_72_11_n_13 | mul_72_11_n_331) & (mul_72_11_n_249 | mul_72_11_n_343));
 assign mul_72_11_n_610 = ~((mul_72_11_n_13 | mul_72_11_n_370) & (mul_72_11_n_249 | mul_72_11_n_371));
 assign mul_72_11_n_609 = ~((mul_72_11_n_13 | mul_72_11_n_175) & (mul_72_11_n_249 | mul_72_11_n_150));
 assign mul_72_11_n_608 = ~((mul_72_11_n_13 | mul_72_11_n_356) & (mul_72_11_n_249 | mul_72_11_n_355));
 assign mul_72_11_n_607 = ~((mul_72_11_n_13 | mul_72_11_n_200) & (mul_72_11_n_249 | mul_72_11_n_199));
 assign mul_72_11_n_606 = ~((mul_72_11_n_13 | mul_72_11_n_332) & (mul_72_11_n_249 | mul_72_11_n_331));
 assign mul_72_11_n_605 = ~((mul_72_11_n_412 | mul_72_11_n_152) & (mul_72_11_n_255 | mul_72_11_n_151));
 assign mul_72_11_n_604 = ~((mul_72_11_n_13 | mul_72_11_n_218) & (mul_72_11_n_249 | mul_72_11_n_217));
 assign mul_72_11_n_603 = ~((mul_72_11_n_412 | mul_72_11_n_347) & (mul_72_11_n_255 | mul_72_11_n_278));
 assign mul_72_11_n_602 = ~((mul_72_11_n_411 | mul_72_11_n_375) & (mul_72_11_n_251 | mul_72_11_n_374));
 assign mul_72_11_n_601 = ~((mul_72_11_n_411 | mul_72_11_n_326) & (mul_72_11_n_251 | mul_72_11_n_340));
 assign mul_72_11_n_600 = ~((mul_72_11_n_411 | mul_72_11_n_104) & (mul_72_11_n_251 | mul_72_11_n_375));
 assign mul_72_11_n_599 = ~((mul_72_11_n_411 | mul_72_11_n_312) & (mul_72_11_n_251 | mul_72_11_n_327));
 assign mul_72_11_n_598 = ~((mul_72_11_n_411 | mul_72_11_n_100) & (mul_72_11_n_251 | mul_72_11_n_104));
 assign mul_72_11_n_597 = ~((mul_72_11_n_411 | mul_72_11_n_340) & (mul_72_11_n_251 | mul_72_11_n_339));
 assign mul_72_11_n_596 = ~((mul_72_11_n_411 | mul_72_11_n_202) & (mul_72_11_n_251 | mul_72_11_n_100));
 assign mul_72_11_n_595 = ~((mul_72_11_n_411 | mul_72_11_n_311) & (mul_72_11_n_251 | mul_72_11_n_312));
 assign mul_72_11_n_594 = ~((mul_72_11_n_411 | mul_72_11_n_293) & (mul_72_11_n_251 | mul_72_11_n_311));
 assign mul_72_11_n_593 = ~((mul_72_11_n_411 | mul_72_11_n_184) & (mul_72_11_n_251 | mul_72_11_n_204));
 assign mul_72_11_n_592 = ~((mul_72_11_n_411 | mul_72_11_n_351) & (mul_72_11_n_251 | mul_72_11_n_352));
 assign mul_72_11_n_591 = ~((mul_72_11_n_411 | mul_72_11_n_163) & (mul_72_11_n_251 | mul_72_11_n_164));
 assign mul_72_11_n_590 = ~((mul_72_11_n_411 | mul_72_11_n_164) & (mul_72_11_n_251 | mul_72_11_n_183));
 assign mul_72_11_n_589 = ~((mul_72_11_n_411 | mul_72_11_n_183) & (mul_72_11_n_251 | mul_72_11_n_184));
 assign mul_72_11_n_588 = ~((mul_72_11_n_411 | mul_72_11_n_204) & (mul_72_11_n_251 | mul_72_11_n_202));
 assign mul_72_11_n_587 = ~((mul_72_11_n_411 | mul_72_11_n_339) & (mul_72_11_n_251 | mul_72_11_n_351));
 assign mul_72_11_n_586 = ~((mul_72_11_n_411 | mul_72_11_n_149) & (mul_72_11_n_251 | mul_72_11_n_163));
 assign mul_72_11_n_585 = ~((mul_72_11_n_412 | mul_72_11_n_319) & (mul_72_11_n_255 | mul_72_11_n_347));
 assign mul_72_11_n_584 = ~((mul_72_11_n_13 | mul_72_11_n_179) & (mul_72_11_n_249 | mul_72_11_n_200));
 assign mul_72_11_n_583 = ~((mul_72_11_n_13 | mul_72_11_n_355) & (mul_72_11_n_249 | mul_72_11_n_370));
 assign mul_72_11_n_582 = ~((mul_72_11_n_13 | mul_72_11_n_316) & (mul_72_11_n_249 | mul_72_11_n_332));
 assign mul_72_11_n_581 = ~((mul_72_11_n_412 | mul_72_11_n_135) & (mul_72_11_n_255 | mul_72_11_n_152));
 assign mul_72_11_n_580 = ~((mul_72_11_n_13 | mul_72_11_n_344) & (mul_72_11_n_249 | mul_72_11_n_356));
 assign mul_72_11_n_579 = ~((mul_72_11_n_13 | mul_72_11_n_300) & (mul_72_11_n_249 | mul_72_11_n_315));
 assign mul_72_11_n_578 = ~((mul_72_11_n_412 | mul_72_11_n_134) & (mul_72_11_n_255 | mul_72_11_n_135));
 assign mul_72_11_n_577 = ~((mul_72_11_n_412 | mul_72_11_n_83) & (mul_72_11_n_255 | mul_72_11_n_319));
 assign mul_72_11_n_576 = ~((mul_72_11_n_412 | mul_72_11_n_303) & (mul_72_11_n_255 | mul_72_11_n_302));
 assign mul_72_11_n_575 = ~((mul_72_11_n_412 | mul_72_11_n_171) & (mul_72_11_n_255 | mul_72_11_n_172));
 assign mul_72_11_n_574 = ~((mul_72_11_n_412 | mul_72_11_n_219) & (mul_72_11_n_255 | mul_72_11_n_83));
 assign mul_72_11_n_573 = ~((mul_72_11_n_13 | mul_72_11_n_180) & (mul_72_11_n_249 | mul_72_11_n_179));
 assign mul_72_11_n_572 = ~((mul_72_11_n_13 | mul_72_11_n_291) & (mul_72_11_n_249 | mul_72_11_n_284));
 assign mul_72_11_n_571 = ~((mul_72_11_n_412 | mul_72_11_n_151) & (mul_72_11_n_255 | mul_72_11_n_171));
 assign mul_72_11_n_570 = ~((mul_72_11_n_412 | mul_72_11_n_82) & (mul_72_11_n_255 | mul_72_11_n_121));
 assign mul_72_11_n_569 = ~((mul_72_11_n_412 | mul_72_11_n_278) & (mul_72_11_n_255 | mul_72_11_n_279));
 assign mul_72_11_n_568 = ~((mul_72_11_n_13 | mul_72_11_n_150) & (mul_72_11_n_249 | mul_72_11_n_360));
 assign mul_72_11_n_567 = ~((mul_72_11_n_411 | mul_72_11_n_68) & (mul_72_11_n_251 | mul_72_11_n_149));
 assign mul_72_11_n_566 = ~((mul_72_11_n_411 | mul_72_11_n_352) & (mul_72_11_n_251 | mul_72_11_n_366));
 assign mul_72_11_n_565 = ~((mul_72_11_n_13 | mul_72_11_n_199) & (mul_72_11_n_249 | mul_72_11_n_218));
 assign mul_72_11_n_564 = ~((mul_72_11_n_13 | mul_72_11_n_217) & (mul_72_11_n_249 | mul_72_11_n_175));
 assign mul_72_11_n_563 = ~((mul_72_11_n_411 | mul_72_11_n_277) & (mul_72_11_n_251 | mul_72_11_n_294));
 assign mul_72_11_n_562 = ~((mul_72_11_n_411 | mul_72_11_n_276) & (mul_72_11_n_251 | mul_72_11_n_277));
 assign mul_72_11_n_561 = ~((mul_72_11_n_411 | mul_72_11_n_294) & (mul_72_11_n_251 | mul_72_11_n_293));
 assign mul_72_11_n_560 = ~((mul_72_11_n_411 | mul_72_11_n_327) & (mul_72_11_n_251 | mul_72_11_n_326));
 assign mul_72_11_n_555 = ~((mul_72_11_n_411 | mul_72_11_n_374) & (mul_72_11_n_251 | mul_72_11_n_276));
 assign mul_72_11_n_553 = ~((mul_72_11_n_391 | mul_72_11_n_147) & (mul_72_11_n_260 | mul_72_11_n_76));
 assign mul_72_11_n_552 = ~((mul_72_11_n_387 | mul_72_11_n_168) & (mul_72_11_n_187 | mul_72_11_n_46));
 assign mul_72_11_n_551 = ~((mul_72_11_n_10 | mul_72_11_n_297) & (mul_72_11_n_250 | mul_72_11_n_244));
 assign mul_72_11_n_550 = ~((mul_72_11_n_392 | mul_72_11_n_108) & (mul_72_11_n_262 | mul_72_11_n_72));
 assign mul_72_11_n_549 = ~((mul_72_11_n_266 | (mul_72_11_n_223 | mul_72_11_n_0)) & (mul_72_11_n_265
    | mul_72_11_n_230));
 assign mul_72_11_n_547 = ~((mul_72_11_n_387 | mul_72_11_n_318) & (mul_72_11_n_317 | mul_72_11_n_46));
 assign mul_72_11_n_546 = ~((mul_72_11_n_390 | mul_72_11_n_102) & (mul_72_11_n_259 | mul_72_11_n_113));
 assign mul_72_11_n_545 = ~((mul_72_11_n_387 | mul_72_11_n_305) & (mul_72_11_n_306 | mul_72_11_n_46));
 assign mul_72_11_n_544 = ~((mul_72_11_n_387 | mul_72_11_n_304) & (mul_72_11_n_376 | mul_72_11_n_46));
 assign mul_72_11_n_543 = ~((mul_72_11_n_387 | mul_72_11_n_372) & (mul_72_11_n_373 | mul_72_11_n_46));
 assign mul_72_11_n_542 = ~((mul_72_11_n_392 | mul_72_11_n_131) & (mul_72_11_n_262 | mul_72_11_n_120));
 assign mul_72_11_n_541 = ~((mul_72_11_n_387 | mul_72_11_n_334) & (mul_72_11_n_333 | mul_72_11_n_46));
 assign mul_72_11_n_540 = ~((mul_72_11_n_387 | mul_72_11_n_270) & (mul_72_11_n_269 | mul_72_11_n_46));
 assign mul_72_11_n_539 = ~((mul_72_11_n_387 | mul_72_11_n_89) & (mul_72_11_n_95 | mul_72_11_n_46));
 assign mul_72_11_n_538 = ~((mul_72_11_n_392 | mul_72_11_n_120) & (mul_72_11_n_262 | mul_72_11_n_119));
 assign mul_72_11_n_537 = ~((mul_72_11_n_387 | mul_72_11_n_333) & (mul_72_11_n_346 | mul_72_11_n_46));
 assign mul_72_11_n_536 = ~((mul_72_11_n_387 | mul_72_11_n_325) & (mul_72_11_n_159 | mul_72_11_n_46));
 assign mul_72_11_n_535 = ~((mul_72_11_n_387 | mul_72_11_n_288) & (mul_72_11_n_287 | mul_72_11_n_46));
 assign mul_72_11_n_534 = ~((mul_72_11_n_387 | mul_72_11_n_363) & (mul_72_11_n_292 | mul_72_11_n_46));
 assign mul_72_11_n_533 = ~((mul_72_11_n_387 | mul_72_11_n_346) & (mul_72_11_n_345 | mul_72_11_n_46));
 assign mul_72_11_n_532 = ~((mul_72_11_n_387 | mul_72_11_n_357) & (mul_72_11_n_358 | mul_72_11_n_46));
 assign mul_72_11_n_531 = ~((mul_72_11_n_387 | mul_72_11_n_187) & (mul_72_11_n_188 | mul_72_11_n_46));
 assign mul_72_11_n_530 = ~((mul_72_11_n_390 | mul_72_11_n_94) & (mul_72_11_n_259 | mul_72_11_n_101));
 assign mul_72_11_n_529 = ~((mul_72_11_n_387 | mul_72_11_n_207) & (mul_72_11_n_206 | mul_72_11_n_46));
 assign mul_72_11_n_528 = ~((mul_72_11_n_387 | mul_72_11_n_362) & (mul_72_11_n_304 | mul_72_11_n_46));
 assign mul_72_11_n_527 = ~((mul_72_11_n_387 | mul_72_11_n_373) & (mul_72_11_n_363 | mul_72_11_n_46));
 assign mul_72_11_n_526 = ~((mul_72_11_n_10 | mul_72_11_n_368) & (mul_72_11_n_250 | mul_72_11_n_297));
 assign mul_72_11_n_525 = ~((mul_72_11_n_387 | mul_72_11_n_287) & (mul_72_11_n_305 | mul_72_11_n_46));
 assign mul_72_11_n_524 = ~((mul_72_11_n_387 | mul_72_11_n_292) & (mul_72_11_n_362 | mul_72_11_n_46));
 assign mul_72_11_n_523 = ~((mul_72_11_n_387 | mul_72_11_n_206) & (mul_72_11_n_89 | mul_72_11_n_46));
 assign mul_72_11_n_522 = ~((mul_72_11_n_392 | mul_72_11_n_119) & (mul_72_11_n_262 | mul_72_11_n_108));
 assign mul_72_11_n_521 = ~((mul_72_11_n_387 | mul_72_11_n_95) & (mul_72_11_n_325 | mul_72_11_n_46));
 assign mul_72_11_n_520 = ~((mul_72_11_n_387 | mul_72_11_n_188) & (mul_72_11_n_207 | mul_72_11_n_46));
 assign mul_72_11_n_519 = ~((mul_72_11_n_392 | mul_72_11_n_139) & (mul_72_11_n_262 | mul_72_11_n_130));
 assign mul_72_11_n_518 = ~((mul_72_11_n_387 | mul_72_11_n_159) & (mul_72_11_n_270 | mul_72_11_n_46));
 assign mul_72_11_n_517 = ~((mul_72_11_n_392 | mul_72_11_n_130) & (mul_72_11_n_262 | mul_72_11_n_131));
 assign mul_72_11_n_516 = ~((mul_72_11_n_392 | mul_72_11_n_236) & (mul_72_11_n_262 | mul_72_11_n_139));
 assign mul_72_11_n_515 = ~((mul_72_11_n_391 | mul_72_11_n_112) & (mul_72_11_n_260 | mul_72_11_n_123));
 assign mul_72_11_n_514 = ~((mul_72_11_n_391 | mul_72_11_n_122) & (mul_72_11_n_260 | mul_72_11_n_147));
 assign mul_72_11_n_513 = ~((mul_72_11_n_391 | mul_72_11_n_123) & (mul_72_11_n_260 | mul_72_11_n_122));
 assign mul_72_11_n_512 = ~((mul_72_11_n_391 | mul_72_11_n_87) & (mul_72_11_n_260 | mul_72_11_n_96));
 assign mul_72_11_n_511 = ~((mul_72_11_n_391 | mul_72_11_n_80) & (mul_72_11_n_260 | mul_72_11_n_86));
 assign mul_72_11_n_510 = ~((mul_72_11_n_387 | mul_72_11_n_345) & (mul_72_11_n_357 | mul_72_11_n_46));
 assign mul_72_11_n_509 = ~((mul_72_11_n_391 | mul_72_11_n_111) & (mul_72_11_n_260 | mul_72_11_n_112));
 assign mul_72_11_n_508 = ~((mul_72_11_n_391 | mul_72_11_n_97) & (mul_72_11_n_260 | mul_72_11_n_111));
 assign mul_72_11_n_507 = ~((mul_72_11_n_391 | mul_72_11_n_88) & (mul_72_11_n_260 | mul_72_11_n_87));
 assign mul_72_11_n_506 = ~((mul_72_11_n_391 | mul_72_11_n_86) & (mul_72_11_n_260 | mul_72_11_n_88));
 assign mul_72_11_n_505 = ~((mul_72_11_n_391 | mul_72_11_n_96) & (mul_72_11_n_260 | mul_72_11_n_97));
 assign mul_72_11_n_504 = ~((mul_72_11_n_387 | mul_72_11_n_306) & (mul_72_11_n_318 | mul_72_11_n_46));
 assign mul_72_11_n_503 = ~((mul_72_11_n_390 | mul_72_11_n_129) & (mul_72_11_n_259 | mul_72_11_n_143));
 assign mul_72_11_n_502 = ~((mul_72_11_n_390 | mul_72_11_n_166) & (mul_72_11_n_259 | mul_72_11_n_201));
 assign mul_72_11_n_501 = ~((mul_72_11_n_387 | mul_72_11_n_358) & (mul_72_11_n_372 | mul_72_11_n_46));
 assign mul_72_11_n_500 = ~((mul_72_11_n_390 | mul_72_11_n_101) & (mul_72_11_n_259 | mul_72_11_n_102));
 assign mul_72_11_n_499 = ~((mul_72_11_n_387 | mul_72_11_n_269) & (mul_72_11_n_288 | mul_72_11_n_46));
 assign mul_72_11_n_498 = ~((mul_72_11_n_390 | mul_72_11_n_143) & (mul_72_11_n_259 | mul_72_11_n_142));
 assign mul_72_11_n_497 = ~((mul_72_11_n_390 | mul_72_11_n_77) & (mul_72_11_n_259 | mul_72_11_n_94));
 assign mul_72_11_n_496 = ~((mul_72_11_n_390 | mul_72_11_n_113) & (mul_72_11_n_259 | mul_72_11_n_114));
 assign mul_72_11_n_495 = ~((mul_72_11_n_390 | mul_72_11_n_114) & (mul_72_11_n_259 | mul_72_11_n_128));
 assign mul_72_11_n_494 = ~((mul_72_11_n_390 | mul_72_11_n_128) & (mul_72_11_n_259 | mul_72_11_n_129));
 assign mul_72_11_n_493 = ~((mul_72_11_n_390 | mul_72_11_n_142) & (mul_72_11_n_259 | mul_72_11_n_165));
 assign mul_72_11_n_492 = ~((mul_72_11_n_390 | mul_72_11_n_165) & (mul_72_11_n_259 | mul_72_11_n_166));
 assign mul_72_11_n_491 = ~((mul_72_11_n_11 | mul_72_11_n_321) & (mul_72_11_n_254 | mul_72_11_n_336));
 assign mul_72_11_n_490 = ~((mul_72_11_n_11 | mul_72_11_n_110) & (mul_72_11_n_254 | mul_72_11_n_107));
 assign mul_72_11_n_489 = ~((mul_72_11_n_387 | mul_72_11_n_317) & (mul_72_11_n_334 | mul_72_11_n_46));
 assign mul_72_11_n_488 = ~((mul_72_11_n_388 & mul_72_11_n_348) | (mul_72_11_n_252 & mul_72_11_n_227));
 assign mul_72_11_n_487 = ~((mul_72_11_n_11 | mul_72_11_n_336) & (mul_72_11_n_254 | mul_72_11_n_226));
 assign mul_72_11_n_486 = ~((mul_72_11_n_389 | mul_72_11_n_154) & (mul_72_11_n_253 | mul_72_11_n_169));
 assign mul_72_11_n_485 = ~((mul_72_11_n_10 | mul_72_11_n_329) & (mul_72_11_n_250 | mul_72_11_n_341));
 assign mul_72_11_n_484 = ~((mul_72_11_n_10 | mul_72_11_n_280) & (mul_72_11_n_250 | mul_72_11_n_298));
 assign mul_72_11_n_483 = ~((mul_72_11_n_10 | mul_72_11_n_118) & (mul_72_11_n_250 | mul_72_11_n_273));
 assign mul_72_11_n_482 = ~((mul_72_11_n_389 | mul_72_11_n_203) & (mul_72_11_n_253 | mul_72_11_n_268));
 assign mul_72_11_n_481 = ~((mul_72_11_n_11 | mul_72_11_n_185) & (mul_72_11_n_254 | mul_72_11_n_208));
 assign mul_72_11_n_480 = ~((mul_72_11_n_11 | mul_72_11_n_186) & (mul_72_11_n_254 | mul_72_11_n_185));
 assign mul_72_11_n_479 = ~((mul_72_11_n_11 | mul_72_11_n_158) & (mul_72_11_n_254 | mul_72_11_n_186));
 assign mul_72_11_n_478 = ~((mul_72_11_n_11 | mul_72_11_n_144) & (mul_72_11_n_254 | mul_72_11_n_214));
 assign mul_72_11_n_477 = ~((mul_72_11_n_11 | mul_72_11_n_361) & (mul_72_11_n_254 | mul_72_11_n_286));
 assign mul_72_11_n_476 = ~((mul_72_11_n_11 | mul_72_11_n_214) & (mul_72_11_n_254 | mul_72_11_n_158));
 assign mul_72_11_n_475 = ~((mul_72_11_n_11 | mul_72_11_n_350) & (mul_72_11_n_254 | mul_72_11_n_361));
 assign mul_72_11_n_474 = ~((mul_72_11_n_11 | mul_72_11_n_322) & (mul_72_11_n_254 | mul_72_11_n_321));
 assign mul_72_11_n_473 = ~((mul_72_11_n_11 | mul_72_11_n_145) & (mul_72_11_n_254 | mul_72_11_n_144));
 assign mul_72_11_n_472 = ~((mul_72_11_n_11 | mul_72_11_n_307) & (mul_72_11_n_254 | mul_72_11_n_322));
 assign mul_72_11_n_471 = ~((mul_72_11_n_11 | mul_72_11_n_133) & (mul_72_11_n_254 | mul_72_11_n_145));
 assign mul_72_11_n_470 = ~((mul_72_11_n_11 | mul_72_11_n_107) & (mul_72_11_n_254 | mul_72_11_n_350));
 assign mul_72_11_n_469 = ~((mul_72_11_n_389 | mul_72_11_n_324) & (mul_72_11_n_253 | mul_72_11_n_338));
 assign mul_72_11_n_468 = ~((mul_72_11_n_389 | mul_72_11_n_323) & (mul_72_11_n_253 | mul_72_11_n_324));
 assign mul_72_11_n_467 = ~((mul_72_11_n_389 | mul_72_11_n_268) & (mul_72_11_n_253 | mul_72_11_n_267));
 assign mul_72_11_n_466 = ~((mul_72_11_n_389 | mul_72_11_n_337) & (mul_72_11_n_253 | mul_72_11_n_349));
 assign mul_72_11_n_465 = ~((mul_72_11_n_11 | mul_72_11_n_308) & (mul_72_11_n_254 | mul_72_11_n_307));
 assign mul_72_11_n_464 = ~((mul_72_11_n_389 | mul_72_11_n_309) & (mul_72_11_n_253 | mul_72_11_n_310));
 assign mul_72_11_n_463 = ~((mul_72_11_n_389 | mul_72_11_n_178) & (mul_72_11_n_253 | mul_72_11_n_203));
 assign mul_72_11_n_462 = ~((mul_72_11_n_389 | mul_72_11_n_310) & (mul_72_11_n_253 | mul_72_11_n_323));
 assign mul_72_11_n_461 = ~((mul_72_11_n_389 | mul_72_11_n_215) & (mul_72_11_n_253 | mul_72_11_n_178));
 assign mul_72_11_n_460 = ~((mul_72_11_n_389 | mul_72_11_n_216) & (mul_72_11_n_253 | mul_72_11_n_215));
 assign mul_72_11_n_459 = ~((mul_72_11_n_389 | mul_72_11_n_196) & (mul_72_11_n_253 | mul_72_11_n_216));
 assign mul_72_11_n_458 = ~((mul_72_11_n_389 | mul_72_11_n_170) & (mul_72_11_n_253 | mul_72_11_n_195));
 assign mul_72_11_n_457 = ~((mul_72_11_n_11 | mul_72_11_n_286) & (mul_72_11_n_254 | mul_72_11_n_285));
 assign mul_72_11_n_456 = ~((mul_72_11_n_389 | mul_72_11_n_195) & (mul_72_11_n_253 | mul_72_11_n_196));
 assign mul_72_11_n_455 = ~((mul_72_11_n_11 | mul_72_11_n_285) & (mul_72_11_n_254 | mul_72_11_n_308));
 assign mul_72_11_n_454 = ~((mul_72_11_n_389 | mul_72_11_n_169) & (mul_72_11_n_253 | mul_72_11_n_170));
 assign mul_72_11_n_453 = ~((mul_72_11_n_389 | mul_72_11_n_338) & (mul_72_11_n_253 | mul_72_11_n_337));
 assign mul_72_11_n_452 = ~((mul_72_11_n_389 | mul_72_11_n_69) & (mul_72_11_n_253 | mul_72_11_n_138));
 assign mul_72_11_n_451 = ~((mul_72_11_n_389 | mul_72_11_n_138) & (mul_72_11_n_253 | mul_72_11_n_153));
 assign mul_72_11_n_450 = ~((mul_72_11_n_11 | mul_72_11_n_209) & (mul_72_11_n_254 | mul_72_11_n_110));
 assign mul_72_11_n_449 = ~((mul_72_11_n_389 | mul_72_11_n_289) & (mul_72_11_n_253 | mul_72_11_n_309));
 assign mul_72_11_n_448 = ~((mul_72_11_n_389 | mul_72_11_n_267) & (mul_72_11_n_253 | mul_72_11_n_290));
 assign mul_72_11_n_447 = ~((mul_72_11_n_389 | mul_72_11_n_153) & (mul_72_11_n_253 | mul_72_11_n_154));
 assign mul_72_11_n_446 = ~((mul_72_11_n_10 | mul_72_11_n_354) & (mul_72_11_n_250 | mul_72_11_n_353));
 assign mul_72_11_n_445 = ~((mul_72_11_n_10 | mul_72_11_n_299) & (mul_72_11_n_250 | mul_72_11_n_314));
 assign mul_72_11_n_444 = ~((mul_72_11_n_10 | mul_72_11_n_67) & (mul_72_11_n_250 | mul_72_11_n_157));
 assign mul_72_11_n_443 = ~((mul_72_11_n_10 | mul_72_11_n_342) & (mul_72_11_n_250 | mul_72_11_n_354));
 assign mul_72_11_n_442 = ~((mul_72_11_n_10 | mul_72_11_n_298) & (mul_72_11_n_250 | mul_72_11_n_299));
 assign mul_72_11_n_441 = ~((mul_72_11_n_10 | mul_72_11_n_191) & (mul_72_11_n_250 | mul_72_11_n_192));
 assign mul_72_11_n_440 = ~((mul_72_11_n_11 | mul_72_11_n_70) & (mul_72_11_n_254 | mul_72_11_n_133));
 assign mul_72_11_n_439 = ~((mul_72_11_n_10 | mul_72_11_n_281) & (mul_72_11_n_250 | mul_72_11_n_280));
 assign mul_72_11_n_438 = ~((mul_72_11_n_10 | mul_72_11_n_378) & (mul_72_11_n_250 | mul_72_11_n_281));
 assign mul_72_11_n_437 = ~((mul_72_11_n_10 | mul_72_11_n_341) & (mul_72_11_n_250 | mul_72_11_n_342));
 assign mul_72_11_n_436 = ~((mul_72_11_n_10 | mul_72_11_n_273) & (mul_72_11_n_250 | mul_72_11_n_378));
 assign mul_72_11_n_435 = ~((mul_72_11_n_11 | mul_72_11_n_208) & (mul_72_11_n_254 | mul_72_11_n_209));
 assign mul_72_11_n_434 = ~((mul_72_11_n_389 | mul_72_11_n_290) & (mul_72_11_n_253 | mul_72_11_n_289));
 assign mul_72_11_n_433 = ~((mul_72_11_n_10 | mul_72_11_n_328) & (mul_72_11_n_250 | mul_72_11_n_329));
 assign mul_72_11_n_432 = ~((mul_72_11_n_10 | mul_72_11_n_132) & (mul_72_11_n_250 | mul_72_11_n_118));
 assign mul_72_11_n_431 = ~((mul_72_11_n_10 | mul_72_11_n_213) & (mul_72_11_n_250 | mul_72_11_n_132));
 assign mul_72_11_n_430 = ~((mul_72_11_n_10 | mul_72_11_n_174) & (mul_72_11_n_250 | mul_72_11_n_191));
 assign mul_72_11_n_429 = ~((mul_72_11_n_10 | mul_72_11_n_353) & (mul_72_11_n_250 | mul_72_11_n_369));
 assign mul_72_11_n_428 = ~((mul_72_11_n_10 | mul_72_11_n_313) & (mul_72_11_n_250 | mul_72_11_n_328));
 assign mul_72_11_n_427 = ~((mul_72_11_n_10 | mul_72_11_n_314) & (mul_72_11_n_250 | mul_72_11_n_313));
 assign mul_72_11_n_426 = ~((mul_72_11_n_10 | mul_72_11_n_212) & (mul_72_11_n_250 | mul_72_11_n_213));
 assign mul_72_11_n_425 = ~((mul_72_11_n_10 | mul_72_11_n_192) & (mul_72_11_n_250 | mul_72_11_n_212));
 assign mul_72_11_n_424 = ~((mul_72_11_n_10 | mul_72_11_n_173) & (mul_72_11_n_250 | mul_72_11_n_174));
 assign mul_72_11_n_423 = ~((mul_72_11_n_10 | mul_72_11_n_157) & (mul_72_11_n_250 | mul_72_11_n_173));
 assign mul_72_11_n_422 = ~((mul_72_11_n_10 | mul_72_11_n_369) & (mul_72_11_n_250 | mul_72_11_n_368));
 assign mul_72_11_n_421 = ~mul_72_11_n_420;
 assign mul_72_11_n_419 = ~mul_72_11_n_418;
 assign mul_72_11_n_417 = ~mul_72_11_n_416;
 assign mul_72_11_n_413 = ~mul_72_11_n_414;
 assign mul_72_11_n_410 = ~mul_72_11_n_411;
 assign mul_72_11_n_420 = ~(mul_72_11_n_264 & mul_72_11_n_228);
 assign mul_72_11_n_409 = ~(mul_72_11_n_264 | mul_72_11_n_37);
 assign mul_72_11_n_418 = ~(mul_72_11_n_263 & mul_72_11_n_229);
 assign mul_72_11_n_416 = ~(mul_72_11_n_261 & mul_72_11_n_234);
 assign mul_72_11_n_415 = (mul_72_11_n_398 | mul_72_11_n_238);
 assign mul_72_11_n_414 = (mul_72_11_n_256 | mul_72_11_n_239);
 assign mul_72_11_n_412 = (mul_72_11_n_393 | mul_72_11_n_240);
 assign mul_72_11_n_411 = (mul_72_11_n_394 | mul_72_11_n_243);
 assign mul_72_11_n_407 = ~(mul_72_11_n_249 | mul_72_11_n_37);
 assign mul_72_11_n_406 = ~(mul_72_11_n_251 | mul_72_11_n_37);
 assign mul_72_11_n_405 = ~(mul_72_11_n_257 | mul_72_11_n_37);
 assign mul_72_11_n_404 = ~(mul_72_11_n_255 | mul_72_11_n_37);
 assign mul_72_11_n_403 = ~(mul_72_11_n_399 | mul_72_11_n_37);
 assign mul_72_11_n_401 = ~(mul_72_11_n_263 | mul_72_11_n_37);
 assign mul_72_11_n_400 = ~(mul_72_11_n_261 | mul_72_11_n_37);
 assign mul_72_11_n_399 = ~mul_72_11_n_256;
 assign mul_72_11_n_398 = ~mul_72_11_n_257;
 assign mul_72_11_n_397 = ~mul_72_11_n_261;
 assign mul_72_11_n_396 = ~mul_72_11_n_263;
 assign mul_72_11_n_395 = ~mul_72_11_n_264;
 assign mul_72_11_n_394 = ~mul_72_11_n_251;
 assign mul_72_11_n_393 = ~mul_72_11_n_255;
 assign mul_72_11_n_388 = ~mul_72_11_n_389;
 assign mul_72_11_n_386 = ~mul_72_11_n_387;
 assign mul_72_11_n_385 = ~(mul_72_11_n_265 | mul_72_11_n_37);
 assign mul_72_11_n_392 = ~(mul_72_11_n_262 & mul_72_11_n_233);
 assign mul_72_11_n_391 = ~(mul_72_11_n_260 & mul_72_11_n_235);
 assign mul_72_11_n_390 = (mul_72_11_n_258 | mul_72_11_n_237);
 assign mul_72_11_n_389 = (mul_72_11_n_252 | mul_72_11_n_242);
 assign mul_72_11_n_384 = ~(mul_72_11_n_259 | mul_72_11_n_37);
 assign mul_72_11_n_383 = ~(mul_72_11_n_250 | mul_72_11_n_37);
 assign mul_72_11_n_382 = ~(mul_72_11_n_262 | mul_72_11_n_37);
 assign mul_72_11_n_381 = ~(mul_72_11_n_254 | mul_72_11_n_37);
 assign mul_72_11_n_380 = ~(mul_72_11_n_253 | mul_72_11_n_37);
 assign mul_72_11_n_379 = ~(mul_72_11_n_260 | mul_72_11_n_37);
 assign mul_72_11_n_377 = ~mul_72_11_n_376;
 assign mul_72_11_n_366 = ~mul_72_11_n_365;
 assign mul_72_11_n_349 = ~mul_72_11_n_348;
 assign mul_72_11_n_296 = ~mul_72_11_n_295;
 assign mul_72_11_n_275 = ~mul_72_11_n_274;
 assign mul_72_11_n_266 = ~mul_72_11_n_265;
 assign mul_72_11_n_258 = ~mul_72_11_n_259;
 assign mul_72_11_n_252 = ~mul_72_11_n_253;
 assign mul_72_11_n_235 = ~((mul_72_11_n_47 & ~n_408) | (n_407 & n_408));
 assign mul_72_11_n_234 = ~((mul_72_11_n_24 & ~n_406) | (n_405 & n_406));
 assign mul_72_11_n_233 = ~((mul_72_11_n_49 & ~n_404) | (n_403 & n_404));
 assign mul_72_11_n_229 = ~((mul_72_11_n_28 & ~n_402) | (n_401 & n_402));
 assign mul_72_11_n_228 = ~((mul_72_11_n_55 & ~n_400) | (n_399 & n_400));
 assign mul_72_11_n_223 = ~(n_397 ^ n_398);
 assign mul_72_11_n_265 = ((mul_72_11_n_55 & ~n_398) | (n_399 & n_398));
 assign mul_72_11_n_264 = ~(n_401 ^ n_400);
 assign mul_72_11_n_263 = ~(n_403 ^ n_402);
 assign mul_72_11_n_262 = ~(n_405 ^ n_404);
 assign mul_72_11_n_261 = ~(n_407 ^ n_406);
 assign mul_72_11_n_177 = ~mul_72_11_n_176;
 assign mul_72_11_n_168 = ~mul_72_11_n_167;
 assign mul_72_11_n_106 = ~mul_72_11_n_105;
 assign mul_72_11_n_63 = ~(mul_72_11_n_38 & mul_72_11_n_37);
 assign mul_72_11_n_62 = ~(mul_72_11_n_24 & mul_72_11_n_37);
 assign mul_72_11_n_61 = ~(mul_72_11_n_45 & mul_72_11_n_37);
 assign mul_72_11_n_60 = ~(mul_72_11_n_44 & mul_72_11_n_37);
 assign mul_72_11_n_59 = ~(mul_72_11_n_39 & mul_72_11_n_37);
 assign {out1[0]} = ~(mul_72_11_n_46 | mul_72_11_n_37);
 assign mul_72_11_n_55 = ~n_399;
 assign mul_72_11_n_49 = ~n_403;
 assign mul_72_11_n_47 = ~n_407;
 assign mul_72_11_n_28 = ~n_401;
 assign mul_72_11_n_24 = ~n_405;
 assign mul_72_11_n_15 = ~(~(mul_72_11_n_415 | mul_72_11_n_367) | (mul_72_11_n_398 & mul_72_11_n_232));
 assign mul_72_11_n_14 = ~(~(mul_72_11_n_412 | mul_72_11_n_320) | (mul_72_11_n_393 & mul_72_11_n_224));
 assign mul_72_11_n_13 = ~(mul_72_11_n_249 & ~mul_72_11_n_246);
 assign mul_72_11_n_12 = ~(~(mul_72_11_n_390 | mul_72_11_n_201) | (mul_72_11_n_258 & mul_72_11_n_81));
 assign mul_72_11_n_11 = ~(mul_72_11_n_254 & ~mul_72_11_n_241);
 assign mul_72_11_n_10 = ~(mul_72_11_n_250 & ~mul_72_11_n_245);
 assign mul_72_11_n_3 = ~(mul_72_11_n_49 & ~n_402);
 assign mul_72_11_n_2 = ~(mul_72_11_n_47 & ~n_406);
 assign mul_72_11_n_1 = ~(mul_72_11_n_28 & ~n_400);
 assign n_429 = ~(add_59_2_n_68 ^ add_59_2_n_4);
 assign n_430 = ~(add_59_2_n_58 ^ add_59_2_n_30);
 assign n_431 = ~(add_59_2_n_52 ^ add_59_2_n_36);
 assign n_432 = ~(add_59_2_n_11 ^ add_59_2_n_37);
 assign n_433 = ~(add_59_2_n_42 ^ add_59_2_n_31);
 assign n_434 = ~((add_59_2_n_33 & ~add_59_2_n_16) | (add_59_2_n_5 & add_59_2_n_16));
 assign n_435 = ({in8[0]} ^ {in9[0]});
 assign n_436 = ~(add_63_2_n_68 ^ add_63_2_n_4);
 assign n_437 = ~(add_63_2_n_58 ^ add_63_2_n_30);
 assign n_438 = ~(add_63_2_n_52 ^ add_63_2_n_36);
 assign n_439 = ~(add_63_2_n_11 ^ add_63_2_n_37);
 assign n_440 = ~(add_63_2_n_42 ^ add_63_2_n_31);
 assign n_441 = ~((add_63_2_n_33 & ~add_63_2_n_16) | (add_63_2_n_5 & add_63_2_n_16));
 assign n_442 = ({in5[0]} ^ {in6[0]});
 assign n_443 = (csa_tree_add_69_2_groupi_n_1428 ^ csa_tree_add_69_2_groupi_n_54);
 assign n_444 = (csa_tree_add_69_2_groupi_n_93 ^ csa_tree_add_69_2_groupi_n_52);
 assign n_445 = ~(csa_tree_add_69_2_groupi_n_1303 ^ csa_tree_add_69_2_groupi_n_1361);
 assign n_446 = ~(csa_tree_add_69_2_groupi_n_1255 ^ csa_tree_add_69_2_groupi_n_1219);
 assign n_447 = ((csa_tree_add_69_2_groupi_n_967 & ~csa_tree_add_69_2_groupi_n_1013) | (csa_tree_add_69_2_groupi_n_966
    & csa_tree_add_69_2_groupi_n_1013));
 assign n_448 = ((csa_tree_add_69_2_groupi_n_879 & ~csa_tree_add_69_2_groupi_n_878) | (csa_tree_add_69_2_groupi_n_880
    & csa_tree_add_69_2_groupi_n_878));
 assign n_449 = ~(csa_tree_add_69_2_groupi_n_710 ^ csa_tree_add_69_2_groupi_n_975);
 assign n_450 = (csa_tree_add_69_2_groupi_n_982 ^ csa_tree_add_69_2_groupi_n_714);
 assign n_452 = ~(n_454 & n_451);
 assign n_451 = ~((csa_tree_add_69_2_groupi_n_137 & ~csa_tree_add_69_2_groupi_n_76) | ({in7[0]} & csa_tree_add_69_2_groupi_n_76));
 assign n_454 = ~(csa_tree_add_69_2_groupi_n_427 | n_453);
 assign n_453 = (n_382 ^ csa_tree_add_69_2_groupi_n_80);
 assign n_456 = ~(csa_tree_add_69_2_groupi_n_425 & n_455);
 assign n_455 = ~((csa_tree_add_69_2_groupi_n_162 & ~n_439) | (n_440 & n_439));
 assign n_457 = (n_391 ^ csa_tree_add_69_2_groupi_n_79);
 assign n_458 = ((n_432 & ~csa_tree_add_69_2_groupi_n_128) | (csa_tree_add_69_2_groupi_n_95 & csa_tree_add_69_2_groupi_n_128));
 assign n_459 = ((csa_tree_add_69_2_groupi_n_165 & ~n_429) | (n_430 & n_429));
 assign n_460 = ~((csa_tree_add_69_2_groupi_n_147 & ~csa_tree_add_69_2_groupi_n_75) | ({in4[2]} & csa_tree_add_69_2_groupi_n_75));
 assign n_461 = ~((csa_tree_add_69_2_groupi_n_108 & ~csa_tree_add_69_2_groupi_n_75) | ({in4[1]} & csa_tree_add_69_2_groupi_n_75));
 assign n_462 = (n_441 ^ {in4[6]});
 assign n_463 = ((csa_tree_add_69_2_groupi_n_94 & ~{in7[2]}) | (csa_tree_add_69_2_groupi_n_95 & {in7[2]}));
 assign n_464 = ((n_434 & ~{in7[11]}) | (csa_tree_add_69_2_groupi_n_130 & {in7[11]}));
 assign n_465 = ~((csa_tree_add_69_2_groupi_n_148 & ~n_434) | ({in7[10]} & n_434));
 assign n_466 = ~((csa_tree_add_69_2_groupi_n_140 & ~n_434) | ({in7[8]} & n_434));
 assign n_467 = ((n_434 & ~{in7[7]}) | (csa_tree_add_69_2_groupi_n_130 & {in7[7]}));
 assign n_468 = ~((csa_tree_add_69_2_groupi_n_138 & ~n_434) | ({in7[6]} & n_434));
 assign n_469 = ~((csa_tree_add_69_2_groupi_n_104 & ~n_434) | ({in7[4]} & n_434));
 assign n_470 = ~((csa_tree_add_69_2_groupi_n_106 & ~n_434) | ({in7[5]} & n_434));
 assign n_471 = ((n_434 & ~{in7[2]}) | (csa_tree_add_69_2_groupi_n_130 & {in7[2]}));
 assign n_472 = ((n_434 & ~{in7[1]}) | (csa_tree_add_69_2_groupi_n_130 & {in7[1]}));
 assign n_473 = ((n_432 & ~{in7[3]}) | (csa_tree_add_69_2_groupi_n_95 & {in7[3]}));
 assign n_474 = ((csa_tree_add_69_2_groupi_n_94 & ~{in7[6]}) | (csa_tree_add_69_2_groupi_n_95 & {in7[6]}));
 assign n_475 = ((csa_tree_add_69_2_groupi_n_94 & ~{in7[1]}) | (csa_tree_add_69_2_groupi_n_95 & {in7[1]}));
 assign n_476 = ~((csa_tree_add_69_2_groupi_n_118 & ~csa_tree_add_69_2_groupi_n_75) | ({in4[3]} & csa_tree_add_69_2_groupi_n_75));
 assign n_477 = ((csa_tree_add_69_2_groupi_n_94 & ~{in7[8]}) | (csa_tree_add_69_2_groupi_n_95 & {in7[8]}));
 assign n_478 = ((csa_tree_add_69_2_groupi_n_94 & ~{in7[9]}) | (csa_tree_add_69_2_groupi_n_95 & {in7[9]}));
 assign n_479 = ((csa_tree_add_69_2_groupi_n_75 & ~{in4[11]}) | (csa_tree_add_69_2_groupi_n_131 & {in4[11]}));
 assign n_480 = ((csa_tree_add_69_2_groupi_n_75 & ~csa_tree_add_69_2_groupi_n_123) | (csa_tree_add_69_2_groupi_n_131
    & csa_tree_add_69_2_groupi_n_123));
 assign n_481 = ((csa_tree_add_69_2_groupi_n_94 & ~{in7[5]}) | (csa_tree_add_69_2_groupi_n_95 & {in7[5]}));
 assign n_482 = ((csa_tree_add_69_2_groupi_n_94 & ~{in7[7]}) | (csa_tree_add_69_2_groupi_n_95 & {in7[7]}));
 assign n_483 = ~((csa_tree_add_69_2_groupi_n_139 & ~csa_tree_add_69_2_groupi_n_75) | ({in4[8]} & csa_tree_add_69_2_groupi_n_75));
 assign n_484 = (csa_tree_add_69_2_groupi_n_150 ^ csa_tree_add_69_2_groupi_n_75);
 assign n_485 = ((csa_tree_add_69_2_groupi_n_77 & ~csa_tree_add_69_2_groupi_n_165) | (n_382 & csa_tree_add_69_2_groupi_n_165));
 assign n_486 = ((csa_tree_add_69_2_groupi_n_74 & ~n_391) | (csa_tree_add_69_2_groupi_n_73 & n_391));
 assign n_487 = (csa_tree_add_69_2_groupi_n_65 ^ csa_tree_add_69_2_groupi_n_134);
 assign n_488 = ((csa_tree_add_69_2_groupi_n_130 & ~n_433) | (n_434 & n_433));
 assign n_489 = ~(csa_tree_add_69_2_groupi_n_100 ^ csa_tree_add_69_2_groupi_n_75);
 assign n_490 = ((csa_tree_add_69_2_groupi_n_71 & ~n_441) | (n_442 & n_441));
 assign n_491 = ((csa_tree_add_69_2_groupi_n_133 & ~{in4[8]}) | (csa_tree_add_69_2_groupi_n_134 & {in4[8]}));
 assign n_492 = ~((csa_tree_add_69_2_groupi_n_123 & ~csa_tree_add_69_2_groupi_n_133) | ({in4[7]} & csa_tree_add_69_2_groupi_n_133));
 assign n_493 = ~((csa_tree_add_69_2_groupi_n_150 & ~csa_tree_add_69_2_groupi_n_133) | ({in4[4]} & csa_tree_add_69_2_groupi_n_133));
 assign n_494 = ~((csa_tree_add_69_2_groupi_n_105 & ~csa_tree_add_69_2_groupi_n_133) | ({in4[5]} & csa_tree_add_69_2_groupi_n_133));
 assign n_495 = ((csa_tree_add_69_2_groupi_n_67 & ~csa_tree_add_69_2_groupi_n_105) | (csa_tree_add_69_2_groupi_n_66
    & csa_tree_add_69_2_groupi_n_105));
 assign n_496 = ~((csa_tree_add_69_2_groupi_n_104 & ~csa_tree_add_69_2_groupi_n_76) | ({in7[4]} & csa_tree_add_69_2_groupi_n_76));
 assign n_497 = ~((csa_tree_add_69_2_groupi_n_108 & ~csa_tree_add_69_2_groupi_n_67) | ({in4[1]} & csa_tree_add_69_2_groupi_n_67));
 assign n_498 = ~(csa_tree_add_69_2_groupi_n_139 ^ csa_tree_add_69_2_groupi_n_67);
 assign n_499 = (n_382 ^ csa_tree_add_69_2_groupi_n_117);
 assign n_500 = ~((csa_tree_add_69_2_groupi_n_141 & ~csa_tree_add_69_2_groupi_n_76) | ({in7[3]} & csa_tree_add_69_2_groupi_n_76));
 assign n_501 = ~(csa_tree_add_69_2_groupi_n_123 ^ csa_tree_add_69_2_groupi_n_67);
 assign n_502 = ~((csa_tree_add_69_2_groupi_n_150 & ~n_391) | ({in4[4]} & n_391));
 assign n_503 = ((csa_tree_add_69_2_groupi_n_76 & ~csa_tree_add_69_2_groupi_n_138) | (csa_tree_add_69_2_groupi_n_77
    & csa_tree_add_69_2_groupi_n_138));
 assign n_504 = ~((csa_tree_add_69_2_groupi_n_147 & ~n_436) | ({in4[2]} & n_436));
 assign n_505 = ((csa_tree_add_69_2_groupi_n_70 & ~{in7[3]}) | (csa_tree_add_69_2_groupi_n_99 & {in7[3]}));
 assign n_506 = ((n_436 & ~{in4[1]}) | (csa_tree_add_69_2_groupi_n_96 & {in4[1]}));
 assign n_507 = ((csa_tree_add_69_2_groupi_n_70 & ~{in7[5]}) | (csa_tree_add_69_2_groupi_n_64 & {in7[5]}));
 assign n_508 = ~((csa_tree_add_69_2_groupi_n_118 & ~csa_tree_add_69_2_groupi_n_68) | ({in4[3]} & csa_tree_add_69_2_groupi_n_68));
 assign n_509 = ((csa_tree_add_69_2_groupi_n_70 & ~csa_tree_add_69_2_groupi_n_146) | (csa_tree_add_69_2_groupi_n_99
    & csa_tree_add_69_2_groupi_n_146));
 assign n_510 = ~((csa_tree_add_69_2_groupi_n_150 & ~csa_tree_add_69_2_groupi_n_69) | ({in4[4]} & csa_tree_add_69_2_groupi_n_69));
 assign n_511 = ((csa_tree_add_69_2_groupi_n_70 & ~{in7[2]}) | (csa_tree_add_69_2_groupi_n_99 & {in7[2]}));
 assign n_512 = ((csa_tree_add_69_2_groupi_n_147 & ~n_439) | ({in4[2]} & n_439));
 assign n_513 = ((csa_tree_add_69_2_groupi_n_133 & ~{in4[6]}) | (csa_tree_add_69_2_groupi_n_134 & {in4[6]}));
endmodule
