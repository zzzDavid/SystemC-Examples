`timescale 1ps / 1ps
module dut_Mul3Add2u8u8Add3u8u8u8Add3u8u8u8_4(
          in8,
          in7,
          in6,
          in5,
          in4,
          in3,
          in2,
          in1,
          out1,
          clk
);
   input [7:0] in8;
   input [7:0] in7;
   input [7:0] in6;
   input [7:0] in5;
   input [7:0] in4;
   input [7:0] in3;
   input [7:0] in2;
   input [7:0] in1;
   output [28:0] out1;
   input clk;
wire add_51_2_n_0, add_51_2_n_1, add_51_2_n_2, add_51_2_n_3, add_51_2_n_4,
     add_51_2_n_5, add_51_2_n_6, add_51_2_n_7, add_51_2_n_8, add_51_2_n_9,
     add_51_2_n_10, add_51_2_n_11, add_51_2_n_12, add_51_2_n_13, add_51_2_n_14,
     add_51_2_n_15, add_51_2_n_16, add_51_2_n_17, add_51_2_n_18, add_51_2_n_19,
     add_51_2_n_20, add_51_2_n_21, add_51_2_n_24, add_51_2_n_26, add_51_2_n_28,
     add_51_2_n_29, add_51_2_n_31, add_51_2_n_32, add_51_2_n_34, add_51_2_n_35,
     add_51_2_n_36, add_51_2_n_40, csa_tree_add_58_2_groupi_n_0,
     csa_tree_add_58_2_groupi_n_1, csa_tree_add_58_2_groupi_n_2,
     csa_tree_add_58_2_groupi_n_3, csa_tree_add_58_2_groupi_n_4,
     csa_tree_add_58_2_groupi_n_6, csa_tree_add_58_2_groupi_n_7,
     csa_tree_add_58_2_groupi_n_8, csa_tree_add_58_2_groupi_n_9,
     csa_tree_add_58_2_groupi_n_10, csa_tree_add_58_2_groupi_n_11,
     csa_tree_add_58_2_groupi_n_12, csa_tree_add_58_2_groupi_n_13,
     csa_tree_add_58_2_groupi_n_14, csa_tree_add_58_2_groupi_n_15,
     csa_tree_add_58_2_groupi_n_16, csa_tree_add_58_2_groupi_n_18,
     csa_tree_add_58_2_groupi_n_20, csa_tree_add_58_2_groupi_n_22,
     csa_tree_add_58_2_groupi_n_24, csa_tree_add_58_2_groupi_n_26,
     csa_tree_add_58_2_groupi_n_28, csa_tree_add_65_2_groupi_n_0,
     csa_tree_add_65_2_groupi_n_1, csa_tree_add_65_2_groupi_n_2,
     csa_tree_add_65_2_groupi_n_3, csa_tree_add_65_2_groupi_n_4,
     csa_tree_add_65_2_groupi_n_6, csa_tree_add_65_2_groupi_n_7,
     csa_tree_add_65_2_groupi_n_8, csa_tree_add_65_2_groupi_n_9,
     csa_tree_add_65_2_groupi_n_10, csa_tree_add_65_2_groupi_n_11,
     csa_tree_add_65_2_groupi_n_12, csa_tree_add_65_2_groupi_n_13,
     csa_tree_add_65_2_groupi_n_14, csa_tree_add_65_2_groupi_n_15,
     csa_tree_add_65_2_groupi_n_16, csa_tree_add_65_2_groupi_n_18,
     csa_tree_add_65_2_groupi_n_20, csa_tree_add_65_2_groupi_n_22,
     csa_tree_add_65_2_groupi_n_24, csa_tree_add_65_2_groupi_n_26,
     csa_tree_add_65_2_groupi_n_28, mul_68_11_n_0, mul_68_11_n_1, mul_68_11_n_2,
     mul_68_11_n_3, mul_68_11_n_4, mul_68_11_n_5, mul_68_11_n_6, mul_68_11_n_7,
     mul_68_11_n_8, mul_68_11_n_9, mul_68_11_n_10, mul_68_11_n_11,
     mul_68_11_n_12, mul_68_11_n_13, mul_68_11_n_14, mul_68_11_n_15,
     mul_68_11_n_16, mul_68_11_n_17, mul_68_11_n_18, mul_68_11_n_19,
     mul_68_11_n_20, mul_68_11_n_21, mul_68_11_n_22, mul_68_11_n_23,
     mul_68_11_n_24, mul_68_11_n_25, mul_68_11_n_26, mul_68_11_n_27,
     mul_68_11_n_28, mul_68_11_n_29, mul_68_11_n_30, mul_68_11_n_32,
     mul_68_11_n_33, mul_68_11_n_34, mul_68_11_n_35, mul_68_11_n_36,
     mul_68_11_n_37, mul_68_11_n_38, mul_68_11_n_39, mul_68_11_n_40,
     mul_68_11_n_41, mul_68_11_n_42, mul_68_11_n_43, mul_68_11_n_44,
     mul_68_11_n_45, mul_68_11_n_46, mul_68_11_n_47, mul_68_11_n_48,
     mul_68_11_n_49, mul_68_11_n_50, mul_68_11_n_51, mul_68_11_n_52,
     mul_68_11_n_53, mul_68_11_n_54, mul_68_11_n_55, mul_68_11_n_56,
     mul_68_11_n_57, mul_68_11_n_58, mul_68_11_n_59, mul_68_11_n_60,
     mul_68_11_n_61, mul_68_11_n_62, mul_68_11_n_63, mul_68_11_n_64,
     mul_68_11_n_65, mul_68_11_n_66, mul_68_11_n_67, mul_68_11_n_68,
     mul_68_11_n_69, mul_68_11_n_70, mul_68_11_n_71, mul_68_11_n_72,
     mul_68_11_n_73, mul_68_11_n_74, mul_68_11_n_75, mul_68_11_n_76,
     mul_68_11_n_77, mul_68_11_n_78, mul_68_11_n_79, mul_68_11_n_80,
     mul_68_11_n_81, mul_68_11_n_82, mul_68_11_n_83, mul_68_11_n_84,
     mul_68_11_n_85, mul_68_11_n_86, mul_68_11_n_87, mul_68_11_n_88,
     mul_68_11_n_89, mul_68_11_n_90, mul_68_11_n_91, mul_68_11_n_92,
     mul_68_11_n_93, mul_68_11_n_94, mul_68_11_n_95, mul_68_11_n_96,
     mul_68_11_n_97, mul_68_11_n_98, mul_68_11_n_99, mul_68_11_n_100,
     mul_68_11_n_101, mul_68_11_n_102, mul_68_11_n_103, mul_68_11_n_104,
     mul_68_11_n_105, mul_68_11_n_106, mul_68_11_n_107, mul_68_11_n_108,
     mul_68_11_n_109, mul_68_11_n_110, mul_68_11_n_111, mul_68_11_n_112,
     mul_68_11_n_113, mul_68_11_n_114, mul_68_11_n_115, mul_68_11_n_116,
     mul_68_11_n_117, mul_68_11_n_118, mul_68_11_n_119, mul_68_11_n_120,
     mul_68_11_n_121, mul_68_11_n_122, mul_68_11_n_123, mul_68_11_n_124,
     mul_68_11_n_125, mul_68_11_n_126, mul_68_11_n_127, mul_68_11_n_128,
     mul_68_11_n_129, mul_68_11_n_130, mul_68_11_n_131, mul_68_11_n_132,
     mul_68_11_n_133, mul_68_11_n_134, mul_68_11_n_135, mul_68_11_n_136,
     mul_68_11_n_137, mul_68_11_n_138, mul_68_11_n_139, mul_68_11_n_140,
     mul_68_11_n_141, mul_68_11_n_142, mul_68_11_n_143, mul_68_11_n_144,
     mul_68_11_n_145, mul_68_11_n_146, mul_68_11_n_147, mul_68_11_n_148,
     mul_68_11_n_149, mul_68_11_n_150, mul_68_11_n_151, mul_68_11_n_152,
     mul_68_11_n_153, mul_68_11_n_154, mul_68_11_n_155, mul_68_11_n_156,
     mul_68_11_n_157, mul_68_11_n_158, mul_68_11_n_159, mul_68_11_n_160,
     mul_68_11_n_161, mul_68_11_n_162, mul_68_11_n_163, mul_68_11_n_164,
     mul_68_11_n_165, mul_68_11_n_166, mul_68_11_n_167, mul_68_11_n_168,
     mul_68_11_n_169, mul_68_11_n_170, mul_68_11_n_171, mul_68_11_n_172,
     mul_68_11_n_173, mul_68_11_n_174, mul_68_11_n_175, mul_68_11_n_176,
     mul_68_11_n_177, mul_68_11_n_178, mul_68_11_n_179, mul_68_11_n_181,
     mul_68_11_n_182, mul_68_11_n_183, mul_68_11_n_184, mul_68_11_n_185,
     mul_68_11_n_186, mul_68_11_n_187, mul_68_11_n_188, mul_68_11_n_189,
     mul_68_11_n_190, mul_68_11_n_191, mul_68_11_n_192, mul_68_11_n_193,
     mul_68_11_n_194, mul_68_11_n_195, mul_68_11_n_196, mul_68_11_n_197,
     mul_68_11_n_198, mul_68_11_n_199, mul_68_11_n_200, mul_68_11_n_201,
     mul_68_11_n_202, mul_68_11_n_203, mul_68_11_n_204, mul_68_11_n_205,
     mul_68_11_n_206, mul_68_11_n_207, mul_68_11_n_208, mul_68_11_n_209,
     mul_68_11_n_210, mul_68_11_n_211, mul_68_11_n_212, mul_68_11_n_213,
     mul_68_11_n_214, mul_68_11_n_215, mul_68_11_n_216, mul_68_11_n_217,
     mul_68_11_n_220, mul_68_11_n_221, mul_68_11_n_222, mul_68_11_n_223,
     mul_68_11_n_224, mul_68_11_n_225, mul_68_11_n_226, mul_68_11_n_227,
     mul_68_11_n_228, mul_68_11_n_229, mul_68_11_n_230, mul_68_11_n_231,
     mul_68_11_n_232, mul_68_11_n_233, mul_68_11_n_234, mul_68_11_n_235,
     mul_68_11_n_236, mul_68_11_n_237, mul_68_11_n_240, mul_68_11_n_241,
     mul_68_11_n_242, mul_68_11_n_243, mul_68_11_n_244, mul_68_11_n_246,
     mul_68_11_n_248, mul_68_11_n_249, mul_68_11_n_250, mul_68_11_n_251,
     mul_68_11_n_252, mul_68_11_n_253, mul_68_11_n_254, mul_68_11_n_255,
     mul_68_11_n_257, mul_68_11_n_258, mul_68_11_n_259, mul_68_11_n_260,
     mul_68_11_n_261, mul_68_11_n_263, mul_68_11_n_264, mul_68_11_n_265,
     mul_68_11_n_266, mul_68_11_n_267, mul_68_11_n_268, mul_68_11_n_269,
     mul_68_11_n_270, mul_68_11_n_271, mul_68_11_n_272, mul_68_11_n_273,
     mul_68_11_n_274, mul_68_11_n_275, mul_68_11_n_276, mul_68_11_n_277,
     mul_68_11_n_278, mul_68_11_n_279, mul_68_11_n_280, mul_68_11_n_281,
     mul_68_11_n_283, mul_68_11_n_284, mul_68_11_n_285, mul_68_11_n_286,
     mul_68_11_n_287, mul_68_11_n_288, mul_68_11_n_290, mul_68_11_n_291,
     mul_68_11_n_292, mul_68_11_n_293, mul_68_11_n_294, mul_68_11_n_295,
     mul_68_11_n_296, mul_68_11_n_297, mul_68_11_n_298, mul_68_11_n_299,
     mul_68_11_n_301, mul_68_11_n_302, mul_68_11_n_303, mul_68_11_n_304,
     mul_68_11_n_305, mul_68_11_n_306, mul_68_11_n_307, mul_68_11_n_308,
     mul_68_11_n_309, mul_68_11_n_310, mul_68_11_n_311, mul_68_11_n_312,
     mul_68_11_n_313, mul_68_11_n_314, mul_68_11_n_315, mul_68_11_n_316,
     mul_68_11_n_317, mul_68_11_n_318, mul_68_11_n_319, mul_68_11_n_321,
     mul_68_11_n_322, mul_68_11_n_323, mul_68_11_n_324, mul_68_11_n_325,
     mul_68_11_n_326, mul_68_11_n_327, mul_68_11_n_328, mul_68_11_n_329,
     mul_68_11_n_330, mul_68_11_n_331, mul_68_11_n_332, mul_68_11_n_333,
     mul_68_11_n_334, mul_68_11_n_335, mul_68_11_n_336, mul_68_11_n_337,
     mul_68_11_n_340, mul_68_11_n_341, mul_68_11_n_342, mul_68_11_n_343,
     mul_68_11_n_344, mul_68_11_n_346, mul_68_11_n_347, mul_68_11_n_349,
     mul_68_11_n_350, mul_68_11_n_351, mul_68_11_n_352, mul_68_11_n_355,
     mul_68_11_n_357, mul_68_11_n_358, mul_71_11_n_3, mul_71_11_n_4,
     mul_71_11_n_5, mul_71_11_n_6, mul_71_11_n_7, mul_71_11_n_8, mul_71_11_n_9,
     mul_71_11_n_10, mul_71_11_n_11, mul_71_11_n_12, mul_71_11_n_13,
     mul_71_11_n_14, mul_71_11_n_15, mul_71_11_n_16, mul_71_11_n_17,
     mul_71_11_n_18, mul_71_11_n_19, mul_71_11_n_20, mul_71_11_n_21,
     mul_71_11_n_22, mul_71_11_n_23, mul_71_11_n_24, mul_71_11_n_25,
     mul_71_11_n_26, mul_71_11_n_27, mul_71_11_n_28, mul_71_11_n_29,
     mul_71_11_n_30, mul_71_11_n_33, mul_71_11_n_35, mul_71_11_n_36,
     mul_71_11_n_37, mul_71_11_n_38, mul_71_11_n_39, mul_71_11_n_40,
     mul_71_11_n_41, mul_71_11_n_42, mul_71_11_n_43, mul_71_11_n_44,
     mul_71_11_n_45, mul_71_11_n_46, mul_71_11_n_47, mul_71_11_n_48,
     mul_71_11_n_49, mul_71_11_n_50, mul_71_11_n_51, mul_71_11_n_52,
     mul_71_11_n_53, mul_71_11_n_54, mul_71_11_n_55, mul_71_11_n_56,
     mul_71_11_n_57, mul_71_11_n_58, mul_71_11_n_59, mul_71_11_n_60,
     mul_71_11_n_61, mul_71_11_n_62, mul_71_11_n_63, mul_71_11_n_64,
     mul_71_11_n_65, mul_71_11_n_66, mul_71_11_n_67, mul_71_11_n_68,
     mul_71_11_n_69, mul_71_11_n_70, mul_71_11_n_71, mul_71_11_n_72,
     mul_71_11_n_73, mul_71_11_n_74, mul_71_11_n_75, mul_71_11_n_76,
     mul_71_11_n_77, mul_71_11_n_78, mul_71_11_n_79, mul_71_11_n_80,
     mul_71_11_n_81, mul_71_11_n_82, mul_71_11_n_83, mul_71_11_n_84,
     mul_71_11_n_85, mul_71_11_n_86, mul_71_11_n_87, mul_71_11_n_88,
     mul_71_11_n_89, mul_71_11_n_90, mul_71_11_n_91, mul_71_11_n_92,
     mul_71_11_n_93, mul_71_11_n_94, mul_71_11_n_95, mul_71_11_n_96,
     mul_71_11_n_97, mul_71_11_n_98, mul_71_11_n_99, mul_71_11_n_100,
     mul_71_11_n_101, mul_71_11_n_102, mul_71_11_n_103, mul_71_11_n_104,
     mul_71_11_n_105, mul_71_11_n_106, mul_71_11_n_107, mul_71_11_n_108,
     mul_71_11_n_109, mul_71_11_n_110, mul_71_11_n_111, mul_71_11_n_112,
     mul_71_11_n_113, mul_71_11_n_114, mul_71_11_n_115, mul_71_11_n_116,
     mul_71_11_n_117, mul_71_11_n_118, mul_71_11_n_119, mul_71_11_n_120,
     mul_71_11_n_121, mul_71_11_n_122, mul_71_11_n_123, mul_71_11_n_124,
     mul_71_11_n_125, mul_71_11_n_126, mul_71_11_n_127, mul_71_11_n_128,
     mul_71_11_n_129, mul_71_11_n_130, mul_71_11_n_131, mul_71_11_n_132,
     mul_71_11_n_133, mul_71_11_n_134, mul_71_11_n_135, mul_71_11_n_136,
     mul_71_11_n_137, mul_71_11_n_138, mul_71_11_n_139, mul_71_11_n_140,
     mul_71_11_n_141, mul_71_11_n_142, mul_71_11_n_143, mul_71_11_n_144,
     mul_71_11_n_145, mul_71_11_n_146, mul_71_11_n_147, mul_71_11_n_148,
     mul_71_11_n_149, mul_71_11_n_150, mul_71_11_n_151, mul_71_11_n_152,
     mul_71_11_n_153, mul_71_11_n_154, mul_71_11_n_155, mul_71_11_n_156,
     mul_71_11_n_157, mul_71_11_n_158, mul_71_11_n_159, mul_71_11_n_160,
     mul_71_11_n_161, mul_71_11_n_162, mul_71_11_n_163, mul_71_11_n_164,
     mul_71_11_n_165, mul_71_11_n_166, mul_71_11_n_167, mul_71_11_n_168,
     mul_71_11_n_169, mul_71_11_n_170, mul_71_11_n_171, mul_71_11_n_172,
     mul_71_11_n_173, mul_71_11_n_174, mul_71_11_n_175, mul_71_11_n_176,
     mul_71_11_n_177, mul_71_11_n_178, mul_71_11_n_179, mul_71_11_n_180,
     mul_71_11_n_181, mul_71_11_n_182, mul_71_11_n_183, mul_71_11_n_184,
     mul_71_11_n_185, mul_71_11_n_186, mul_71_11_n_187, mul_71_11_n_188,
     mul_71_11_n_189, mul_71_11_n_190, mul_71_11_n_191, mul_71_11_n_192,
     mul_71_11_n_193, mul_71_11_n_194, mul_71_11_n_195, mul_71_11_n_196,
     mul_71_11_n_197, mul_71_11_n_198, mul_71_11_n_199, mul_71_11_n_200,
     mul_71_11_n_201, mul_71_11_n_202, mul_71_11_n_203, mul_71_11_n_204,
     mul_71_11_n_205, mul_71_11_n_206, mul_71_11_n_207, mul_71_11_n_208,
     mul_71_11_n_209, mul_71_11_n_210, mul_71_11_n_211, mul_71_11_n_212,
     mul_71_11_n_213, mul_71_11_n_214, mul_71_11_n_215, mul_71_11_n_216,
     mul_71_11_n_217, mul_71_11_n_218, mul_71_11_n_219, mul_71_11_n_220,
     mul_71_11_n_221, mul_71_11_n_222, mul_71_11_n_223, mul_71_11_n_224,
     mul_71_11_n_225, mul_71_11_n_226, mul_71_11_n_227, mul_71_11_n_228,
     mul_71_11_n_229, mul_71_11_n_230, mul_71_11_n_231, mul_71_11_n_232,
     mul_71_11_n_233, mul_71_11_n_234, mul_71_11_n_235, mul_71_11_n_236,
     mul_71_11_n_237, mul_71_11_n_238, mul_71_11_n_239, mul_71_11_n_240,
     mul_71_11_n_241, mul_71_11_n_242, mul_71_11_n_243, mul_71_11_n_244,
     mul_71_11_n_245, mul_71_11_n_246, mul_71_11_n_247, mul_71_11_n_248,
     mul_71_11_n_249, mul_71_11_n_250, mul_71_11_n_251, mul_71_11_n_252,
     mul_71_11_n_253, mul_71_11_n_255, mul_71_11_n_256, mul_71_11_n_257,
     mul_71_11_n_258, mul_71_11_n_259, mul_71_11_n_260, mul_71_11_n_261,
     mul_71_11_n_262, mul_71_11_n_263, mul_71_11_n_264, mul_71_11_n_265,
     mul_71_11_n_266, mul_71_11_n_267, mul_71_11_n_268, mul_71_11_n_269,
     mul_71_11_n_270, mul_71_11_n_271, mul_71_11_n_272, mul_71_11_n_273,
     mul_71_11_n_274, mul_71_11_n_275, mul_71_11_n_276, mul_71_11_n_277,
     mul_71_11_n_278, mul_71_11_n_279, mul_71_11_n_280, mul_71_11_n_281,
     mul_71_11_n_282, mul_71_11_n_283, mul_71_11_n_284, mul_71_11_n_285,
     mul_71_11_n_286, mul_71_11_n_287, mul_71_11_n_288, mul_71_11_n_289,
     mul_71_11_n_290, mul_71_11_n_291, mul_71_11_n_292, mul_71_11_n_293,
     mul_71_11_n_295, mul_71_11_n_296, mul_71_11_n_297, mul_71_11_n_298,
     mul_71_11_n_299, mul_71_11_n_300, mul_71_11_n_301, mul_71_11_n_302,
     mul_71_11_n_303, mul_71_11_n_304, mul_71_11_n_305, mul_71_11_n_306,
     mul_71_11_n_307, mul_71_11_n_308, mul_71_11_n_309, mul_71_11_n_310,
     mul_71_11_n_311, mul_71_11_n_312, mul_71_11_n_313, mul_71_11_n_314,
     mul_71_11_n_315, mul_71_11_n_316, mul_71_11_n_317, mul_71_11_n_318,
     mul_71_11_n_319, mul_71_11_n_320, mul_71_11_n_321, mul_71_11_n_322,
     mul_71_11_n_323, mul_71_11_n_324, mul_71_11_n_325, mul_71_11_n_326,
     mul_71_11_n_327, mul_71_11_n_328, mul_71_11_n_329, mul_71_11_n_330,
     mul_71_11_n_332, mul_71_11_n_333, mul_71_11_n_334, mul_71_11_n_335,
     mul_71_11_n_336, mul_71_11_n_337, mul_71_11_n_338, mul_71_11_n_339,
     mul_71_11_n_340, mul_71_11_n_341, mul_71_11_n_342, mul_71_11_n_343,
     mul_71_11_n_344, mul_71_11_n_345, mul_71_11_n_346, mul_71_11_n_347,
     mul_71_11_n_348, mul_71_11_n_349, mul_71_11_n_350, mul_71_11_n_351,
     mul_71_11_n_353, mul_71_11_n_354, mul_71_11_n_355, mul_71_11_n_356,
     mul_71_11_n_357, mul_71_11_n_358, mul_71_11_n_359, mul_71_11_n_360,
     mul_71_11_n_361, mul_71_11_n_362, mul_71_11_n_363, mul_71_11_n_364,
     mul_71_11_n_365, mul_71_11_n_366, mul_71_11_n_367, mul_71_11_n_368,
     mul_71_11_n_369, mul_71_11_n_370, mul_71_11_n_371, mul_71_11_n_372,
     mul_71_11_n_373, mul_71_11_n_374, mul_71_11_n_375, mul_71_11_n_376,
     mul_71_11_n_377, mul_71_11_n_379, mul_71_11_n_380, mul_71_11_n_381,
     mul_71_11_n_382, mul_71_11_n_383, mul_71_11_n_384, mul_71_11_n_385,
     mul_71_11_n_386, mul_71_11_n_387, mul_71_11_n_388, mul_71_11_n_389,
     mul_71_11_n_390, mul_71_11_n_391, mul_71_11_n_392, mul_71_11_n_393,
     mul_71_11_n_394, mul_71_11_n_395, mul_71_11_n_396, mul_71_11_n_397,
     mul_71_11_n_398, mul_71_11_n_399, mul_71_11_n_400, mul_71_11_n_401,
     mul_71_11_n_402, mul_71_11_n_403, mul_71_11_n_405, mul_71_11_n_406,
     mul_71_11_n_407, mul_71_11_n_408, mul_71_11_n_409, mul_71_11_n_410,
     mul_71_11_n_411, mul_71_11_n_412, mul_71_11_n_413, mul_71_11_n_414,
     mul_71_11_n_415, mul_71_11_n_416, mul_71_11_n_417, mul_71_11_n_418,
     mul_71_11_n_419, mul_71_11_n_420, mul_71_11_n_421, mul_71_11_n_422,
     mul_71_11_n_423, mul_71_11_n_424, mul_71_11_n_425, mul_71_11_n_426,
     mul_71_11_n_427, mul_71_11_n_428, mul_71_11_n_429, mul_71_11_n_430,
     mul_71_11_n_432, mul_71_11_n_433, mul_71_11_n_434, mul_71_11_n_435,
     mul_71_11_n_436, mul_71_11_n_437, mul_71_11_n_438, mul_71_11_n_439,
     mul_71_11_n_440, mul_71_11_n_441, mul_71_11_n_442, mul_71_11_n_443,
     mul_71_11_n_444, mul_71_11_n_445, mul_71_11_n_446, mul_71_11_n_447,
     mul_71_11_n_448, mul_71_11_n_449, mul_71_11_n_450, mul_71_11_n_451,
     mul_71_11_n_452, mul_71_11_n_453, mul_71_11_n_454, mul_71_11_n_455,
     mul_71_11_n_456, mul_71_11_n_457, mul_71_11_n_458, mul_71_11_n_459,
     mul_71_11_n_460, mul_71_11_n_461, mul_71_11_n_462, mul_71_11_n_463,
     mul_71_11_n_464, mul_71_11_n_465, mul_71_11_n_466, mul_71_11_n_467,
     mul_71_11_n_468, mul_71_11_n_469, mul_71_11_n_470, mul_71_11_n_471,
     mul_71_11_n_472, mul_71_11_n_473, mul_71_11_n_474, mul_71_11_n_475,
     mul_71_11_n_476, mul_71_11_n_477, mul_71_11_n_478, mul_71_11_n_479,
     mul_71_11_n_480, mul_71_11_n_481, mul_71_11_n_483, mul_71_11_n_484,
     mul_71_11_n_485, mul_71_11_n_486, mul_71_11_n_487, mul_71_11_n_488,
     mul_71_11_n_489, mul_71_11_n_490, mul_71_11_n_491, mul_71_11_n_492,
     mul_71_11_n_493, mul_71_11_n_494, mul_71_11_n_495, mul_71_11_n_496,
     mul_71_11_n_498, mul_71_11_n_499, mul_71_11_n_500, mul_71_11_n_501,
     mul_71_11_n_502, mul_71_11_n_504, mul_71_11_n_505, mul_71_11_n_506,
     mul_71_11_n_509, mul_71_11_n_510, mul_71_11_n_511, mul_71_11_n_512,
     mul_71_11_n_515, mul_71_11_n_516, mul_71_11_n_518, mul_71_11_n_519,
     mul_71_11_n_520, mul_71_11_n_522, mul_71_11_n_525, mul_71_11_n_526,
     mul_71_11_n_527, mul_71_11_n_529, mul_71_11_n_530, mul_71_11_n_533,
     mul_71_11_n_534, mul_71_11_n_537, mul_71_11_n_538, mul_71_11_n_541,
     mul_71_11_n_542, n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9, n_10,
     n_11, n_12, n_13, n_14, n_15, n_16, n_17, n_18, n_19, n_20, n_21, n_22,
     n_23, n_24, n_25, clk, n_56, n_57, n_58, n_59, n_60, n_61, n_62, n_63, n_64,
     n_65, n_66, n_67, n_68, n_69, n_70, n_71, n_72, n_73, n_74, n_75, n_76,
     n_77, n_78, n_79, n_144, n_145, n_146, n_147, n_148, n_149, n_150, n_151,
     n_152, n_153, n_154, n_155, n_156, n_157, n_158, n_159, n_160, n_161, n_162,
     n_163, n_164, n_165, n_166, n_167, n_168, n_169, n_170, n_171, n_172, n_173,
     n_174, n_175, n_176, n_177, n_178, n_179, n_180, n_181, n_182, n_183, n_184,
     n_185, n_186, n_187, n_188, n_189, n_190, n_191;
 reg retime_s1_1_reg_reg_N30;
 always @(posedge clk)
         retime_s1_1_reg_reg_N30 <= n_21;
 assign n_56 = retime_s1_1_reg_reg_N30;
 reg retime_s1_2_reg_reg_N30;
 always @(posedge clk)
         retime_s1_2_reg_reg_N30 <= n_168;
 assign n_57 = retime_s1_2_reg_reg_N30;
 reg retime_s1_3_reg_reg_N30;
 always @(posedge clk)
         retime_s1_3_reg_reg_N30 <= n_170;
 assign n_58 = retime_s1_3_reg_reg_N30;
 reg retime_s1_4_reg_reg_N30;
 always @(posedge clk)
         if (mul_68_11_n_333)
         retime_s1_4_reg_reg_N30 <= n_184;
     else
         retime_s1_4_reg_reg_N30 <= mul_68_11_n_351;
 assign mul_71_11_n_24 = retime_s1_4_reg_reg_N30;
 reg retime_s1_5_reg_reg_N30;
 always @(posedge clk)
         retime_s1_5_reg_reg_N30 <= n_179;
 assign n_59 = retime_s1_5_reg_reg_N30;
 reg retime_s1_6_reg_reg_N30;
 always @(posedge clk)
         retime_s1_6_reg_reg_N30 <= n_176;
 assign n_60 = retime_s1_6_reg_reg_N30;
 reg retime_s1_7_reg_reg_N30;
 always @(posedge clk)
         if (mul_68_11_n_322)
         retime_s1_7_reg_reg_N30 <= n_189;
     else
         retime_s1_7_reg_reg_N30 <= mul_68_11_n_311;
 assign mul_71_11_n_29 = retime_s1_7_reg_reg_N30;
 reg retime_s1_8_reg_reg_N30;
 always @(posedge clk)
         if (mul_68_11_n_347)
         retime_s1_8_reg_reg_N30 <= n_183;
     else
         retime_s1_8_reg_reg_N30 <= mul_68_11_n_332;
 assign mul_71_11_n_17 = retime_s1_8_reg_reg_N30;
 reg retime_s1_9_reg_reg_N30;
 always @(posedge clk)
         if (mul_68_11_n_340)
         retime_s1_9_reg_reg_N30 <= n_188;
     else
         retime_s1_9_reg_reg_N30 <= mul_68_11_n_331;
 assign mul_71_11_n_28 = retime_s1_9_reg_reg_N30;
 reg retime_s1_10_reg_reg_N30;
 always @(posedge clk)
         retime_s1_10_reg_reg_N30 <= n_180;
 assign n_61 = retime_s1_10_reg_reg_N30;
 reg retime_s1_11_reg_reg_N30;
 always @(posedge clk)
         if (mul_68_11_n_284)
         retime_s1_11_reg_reg_N30 <= n_186;
     else
         retime_s1_11_reg_reg_N30 <= mul_68_11_n_290;
 assign mul_71_11_n_10 = retime_s1_11_reg_reg_N30;
 reg retime_s1_12_reg_reg_N30;
 always @(posedge clk)
         if (mul_68_11_n_257)
         retime_s1_12_reg_reg_N30 <= n_190;
     else
         retime_s1_12_reg_reg_N30 <= mul_68_11_n_273;
 assign mul_71_11_n_16 = retime_s1_12_reg_reg_N30;
 reg retime_s1_13_reg_reg_N30;
 always @(posedge clk)
         retime_s1_13_reg_reg_N30 <= n_2;
 assign n_62 = retime_s1_13_reg_reg_N30;
 reg retime_s1_14_reg_reg_N30;
 always @(posedge clk)
         retime_s1_14_reg_reg_N30 <= n_166;
 assign n_63 = retime_s1_14_reg_reg_N30;
 reg retime_s1_15_reg_reg_N30;
 always @(posedge clk)
         retime_s1_15_reg_reg_N30 <= n_171;
 assign n_64 = retime_s1_15_reg_reg_N30;
 reg retime_s1_16_reg_reg_N30;
 always @(posedge clk)
         if (mul_68_11_n_237)
         retime_s1_16_reg_reg_N30 <= n_25;
     else
         retime_s1_16_reg_reg_N30 <= mul_68_11_n_255;
 assign mul_71_11_n_14 = retime_s1_16_reg_reg_N30;
 reg retime_s1_17_reg_reg_N30;
 always @(posedge clk)
         if (mul_68_11_n_236)
         retime_s1_17_reg_reg_N30 <= n_0;
     else
         retime_s1_17_reg_reg_N30 <= mul_68_11_n_246;
 assign mul_71_11_n_25 = retime_s1_17_reg_reg_N30;
 reg retime_s1_18_reg_reg_N30;
 always @(posedge clk)
         retime_s1_18_reg_reg_N30 <= n_169;
 assign n_65 = retime_s1_18_reg_reg_N30;
 reg retime_s1_19_reg_reg_N30;
 always @(posedge clk)
         if (mul_68_11_n_318)
         retime_s1_19_reg_reg_N30 <= n_191;
     else
         retime_s1_19_reg_reg_N30 <= mul_68_11_n_292;
 assign mul_71_11_n_8 = retime_s1_19_reg_reg_N30;
 reg retime_s1_20_reg_reg_N30;
 always @(posedge clk)
         retime_s1_20_reg_reg_N30 <= n_24;
 assign n_66 = retime_s1_20_reg_reg_N30;
 reg retime_s1_21_reg_reg_N30;
 always @(posedge clk)
         retime_s1_21_reg_reg_N30 <= n_22;
 assign n_67 = retime_s1_21_reg_reg_N30;
 reg retime_s1_22_reg_reg_N30;
 always @(posedge clk)
         retime_s1_22_reg_reg_N30 <= n_13;
 assign n_68 = retime_s1_22_reg_reg_N30;
 reg retime_s1_23_reg_reg_N30;
 always @(posedge clk)
         retime_s1_23_reg_reg_N30 <= n_177;
 assign mul_71_11_n_22 = retime_s1_23_reg_reg_N30;
 reg retime_s1_24_reg_reg_N30;
 always @(posedge clk)
         retime_s1_24_reg_reg_N30 <= n_1;
 assign n_69 = retime_s1_24_reg_reg_N30;
 reg retime_s1_25_reg_reg_N30;
 always @(posedge clk)
         retime_s1_25_reg_reg_N30 <= n_173;
 assign n_70 = retime_s1_25_reg_reg_N30;
 reg retime_s1_26_reg_reg_N30;
 always @(posedge clk)
         if (mul_68_11_n_350)
         retime_s1_26_reg_reg_N30 <= n_185;
     else
         retime_s1_26_reg_reg_N30 <= mul_68_11_n_319;
 assign mul_71_11_n_26 = retime_s1_26_reg_reg_N30;
 reg retime_s1_27_reg_reg_N30;
 always @(posedge clk)
         retime_s1_27_reg_reg_N30 <= n_172;
 assign n_71 = retime_s1_27_reg_reg_N30;
 reg retime_s1_28_reg_reg_N30;
 always @(posedge clk)
         retime_s1_28_reg_reg_N30 <= n_175;
 assign n_72 = retime_s1_28_reg_reg_N30;
 reg retime_s1_29_reg_reg_N30;
 always @(posedge clk)
         retime_s1_29_reg_reg_N30 <= n_178;
 assign mul_71_11_n_21 = retime_s1_29_reg_reg_N30;
 reg retime_s1_30_reg_reg_N30;
 always @(posedge clk)
         retime_s1_30_reg_reg_N30 <= n_174;
 assign n_73 = retime_s1_30_reg_reg_N30;
 reg retime_s1_31_reg_reg_N30;
 always @(posedge clk)
         if (mul_68_11_n_301)
         retime_s1_31_reg_reg_N30 <= n_187;
     else
         retime_s1_31_reg_reg_N30 <= mul_68_11_n_283;
 assign mul_71_11_n_18 = retime_s1_31_reg_reg_N30;
 assign add_51_2_n_40 = ~(add_51_2_n_8 & (add_51_2_n_34 | add_51_2_n_0));
 assign add_51_2_n_36 = ~(add_51_2_n_5 | (add_51_2_n_32 & (add_51_2_n_16 & add_51_2_n_18)));
 assign add_51_2_n_35 = ~(add_51_2_n_11 & (add_51_2_n_31 | add_51_2_n_7));
 assign add_51_2_n_34 = ~(add_51_2_n_21 | (add_51_2_n_32 & add_51_2_n_16));
 assign add_51_2_n_31 = ~add_51_2_n_32;
 assign add_51_2_n_32 = ~(add_51_2_n_4 & (add_51_2_n_29 | add_51_2_n_12));
 assign add_51_2_n_29 = ~(add_51_2_n_9 | (add_51_2_n_26 & add_51_2_n_2));
 assign add_51_2_n_28 = ~(add_51_2_n_10 & ~(add_51_2_n_26 & add_51_2_n_2));
 assign add_51_2_n_24 = ~(add_51_2_n_21 & add_51_2_n_18);
 assign add_51_2_n_21 = ~(add_51_2_n_3 & (add_51_2_n_1 | add_51_2_n_11));
 assign add_51_2_n_20 = ~(add_51_2_n_7 | ~add_51_2_n_11);
 assign add_51_2_n_19 = ~(add_51_2_n_4 & ~add_51_2_n_12);
 assign add_51_2_n_18 = ~(add_51_2_n_0 | add_51_2_n_6);
 assign add_51_2_n_17 = (add_51_2_n_6 | add_51_2_n_5);
 assign add_51_2_n_16 = ~(add_51_2_n_7 | add_51_2_n_1);
 assign add_51_2_n_15 = ~(add_51_2_n_2 & add_51_2_n_10);
 assign add_51_2_n_14 = ~(add_51_2_n_0 | ~add_51_2_n_8);
 assign add_51_2_n_13 = ~(add_51_2_n_3 & ~add_51_2_n_1);
 assign add_51_2_n_9 = ~add_51_2_n_10;
 assign add_51_2_n_12 = ~({in1[3]} | {in2[3]});
 assign add_51_2_n_11 = ~({in1[4]} & {in2[4]});
 assign add_51_2_n_10 = ~({in1[2]} & {in2[2]});
 assign add_51_2_n_8 = ~({in1[6]} & {in2[6]});
 assign add_51_2_n_7 = ~({in1[4]} | {in2[4]});
 assign add_51_2_n_6 = ~({in1[7]} | {in2[7]});
 assign add_51_2_n_5 = ({in1[7]} & {in2[7]});
 assign add_51_2_n_4 = ~({in1[3]} & {in2[3]});
 assign add_51_2_n_3 = ~({in1[5]} & {in2[5]});
 assign add_51_2_n_2 = ({in1[2]} | {in2[2]});
 assign add_51_2_n_1 = ~({in1[5]} | {in2[5]});
 assign add_51_2_n_0 = ~({in1[6]} | {in2[6]});
 assign n_144 = (csa_tree_add_58_2_groupi_n_28 & csa_tree_add_58_2_groupi_n_14);
 assign n_145 = (csa_tree_add_58_2_groupi_n_28 ^ csa_tree_add_58_2_groupi_n_14);
 assign csa_tree_add_58_2_groupi_n_28 = ((csa_tree_add_58_2_groupi_n_26 & csa_tree_add_58_2_groupi_n_15)
    | ((csa_tree_add_58_2_groupi_n_15 & csa_tree_add_58_2_groupi_n_10) | (csa_tree_add_58_2_groupi_n_10 &
    csa_tree_add_58_2_groupi_n_26)));
 assign n_146 = (csa_tree_add_58_2_groupi_n_15 ^ (csa_tree_add_58_2_groupi_n_10 ^ csa_tree_add_58_2_groupi_n_26));
 assign csa_tree_add_58_2_groupi_n_26 = ((csa_tree_add_58_2_groupi_n_24 & csa_tree_add_58_2_groupi_n_11)
    | ((csa_tree_add_58_2_groupi_n_11 & csa_tree_add_58_2_groupi_n_2) | (csa_tree_add_58_2_groupi_n_2 & csa_tree_add_58_2_groupi_n_24)));
 assign n_147 = (csa_tree_add_58_2_groupi_n_11 ^ (csa_tree_add_58_2_groupi_n_2 ^ csa_tree_add_58_2_groupi_n_24));
 assign csa_tree_add_58_2_groupi_n_24 = ((csa_tree_add_58_2_groupi_n_22 & csa_tree_add_58_2_groupi_n_3)
    | ((csa_tree_add_58_2_groupi_n_3 & csa_tree_add_58_2_groupi_n_12) | (csa_tree_add_58_2_groupi_n_12 &
    csa_tree_add_58_2_groupi_n_22)));
 assign n_148 = (csa_tree_add_58_2_groupi_n_3 ^ (csa_tree_add_58_2_groupi_n_12 ^ csa_tree_add_58_2_groupi_n_22));
 assign csa_tree_add_58_2_groupi_n_22 = ((csa_tree_add_58_2_groupi_n_20 & csa_tree_add_58_2_groupi_n_8)
    | ((csa_tree_add_58_2_groupi_n_8 & csa_tree_add_58_2_groupi_n_13) | (csa_tree_add_58_2_groupi_n_13 &
    csa_tree_add_58_2_groupi_n_20)));
 assign n_149 = (csa_tree_add_58_2_groupi_n_8 ^ (csa_tree_add_58_2_groupi_n_13 ^ csa_tree_add_58_2_groupi_n_20));
 assign csa_tree_add_58_2_groupi_n_20 = ((csa_tree_add_58_2_groupi_n_18 & csa_tree_add_58_2_groupi_n_9)
    | ((csa_tree_add_58_2_groupi_n_9 & csa_tree_add_58_2_groupi_n_6) | (csa_tree_add_58_2_groupi_n_6 & csa_tree_add_58_2_groupi_n_18)));
 assign n_150 = (csa_tree_add_58_2_groupi_n_9 ^ (csa_tree_add_58_2_groupi_n_6 ^ csa_tree_add_58_2_groupi_n_18));
 assign csa_tree_add_58_2_groupi_n_18 = ((csa_tree_add_58_2_groupi_n_16 & csa_tree_add_58_2_groupi_n_7)
    | ((csa_tree_add_58_2_groupi_n_7 & csa_tree_add_58_2_groupi_n_0) | (csa_tree_add_58_2_groupi_n_0 & csa_tree_add_58_2_groupi_n_16)));
 assign n_151 = (csa_tree_add_58_2_groupi_n_7 ^ (csa_tree_add_58_2_groupi_n_0 ^ csa_tree_add_58_2_groupi_n_16));
 assign csa_tree_add_58_2_groupi_n_16 = ((csa_tree_add_58_2_groupi_n_4 & {in5[1]}) | (({in5[1]} & csa_tree_add_58_2_groupi_n_1)
    | (csa_tree_add_58_2_groupi_n_1 & csa_tree_add_58_2_groupi_n_4)));
 assign n_152 = ({in5[1]} ^ (csa_tree_add_58_2_groupi_n_1 ^ csa_tree_add_58_2_groupi_n_4));
 assign csa_tree_add_58_2_groupi_n_14 = (({in4[7]} & {in3[7]}) | (({in3[7]} & {in5[7]}) | ({in5[7]} &
    {in4[7]})));
 assign csa_tree_add_58_2_groupi_n_15 = ({in3[7]} ^ ({in5[7]} ^ {in4[7]}));
 assign csa_tree_add_58_2_groupi_n_12 = (({in4[4]} & {in3[4]}) | (({in3[4]} & {in5[4]}) | ({in5[4]} &
    {in4[4]})));
 assign csa_tree_add_58_2_groupi_n_13 = ({in3[4]} ^ ({in5[4]} ^ {in4[4]}));
 assign csa_tree_add_58_2_groupi_n_10 = (({in4[6]} & {in3[6]}) | (({in3[6]} & {in5[6]}) | ({in5[6]} &
    {in4[6]})));
 assign csa_tree_add_58_2_groupi_n_11 = ({in3[6]} ^ ({in5[6]} ^ {in4[6]}));
 assign csa_tree_add_58_2_groupi_n_8 = (({in4[3]} & {in3[3]}) | (({in3[3]} & {in5[3]}) | ({in5[3]} &
    {in4[3]})));
 assign csa_tree_add_58_2_groupi_n_9 = ({in3[3]} ^ ({in5[3]} ^ {in4[3]}));
 assign csa_tree_add_58_2_groupi_n_6 = (({in4[2]} & {in3[2]}) | (({in3[2]} & {in5[2]}) | ({in5[2]} &
    {in4[2]})));
 assign csa_tree_add_58_2_groupi_n_7 = ({in3[2]} ^ ({in5[2]} ^ {in4[2]}));
 assign csa_tree_add_58_2_groupi_n_4 = (({in3[0]} & {in5[0]}) | (({in5[0]} & {in4[0]}) | ({in4[0]} &
    {in3[0]})));
 assign n_153 = ({in5[0]} ^ ({in4[0]} ^ {in3[0]}));
 assign csa_tree_add_58_2_groupi_n_2 = (({in5[5]} & {in3[5]}) | (({in3[5]} & {in4[5]}) | ({in4[5]} &
    {in5[5]})));
 assign csa_tree_add_58_2_groupi_n_3 = ({in3[5]} ^ ({in4[5]} ^ {in5[5]}));
 assign csa_tree_add_58_2_groupi_n_0 = ({in4[1]} & {in3[1]});
 assign csa_tree_add_58_2_groupi_n_1 = ({in4[1]} ^ {in3[1]});
 assign n_154 = (csa_tree_add_65_2_groupi_n_28 & csa_tree_add_65_2_groupi_n_14);
 assign n_155 = (csa_tree_add_65_2_groupi_n_28 ^ csa_tree_add_65_2_groupi_n_14);
 assign csa_tree_add_65_2_groupi_n_28 = ((csa_tree_add_65_2_groupi_n_26 & csa_tree_add_65_2_groupi_n_10)
    | ((csa_tree_add_65_2_groupi_n_10 & csa_tree_add_65_2_groupi_n_15) | (csa_tree_add_65_2_groupi_n_15 &
    csa_tree_add_65_2_groupi_n_26)));
 assign n_156 = (csa_tree_add_65_2_groupi_n_10 ^ (csa_tree_add_65_2_groupi_n_15 ^ csa_tree_add_65_2_groupi_n_26));
 assign csa_tree_add_65_2_groupi_n_26 = ((csa_tree_add_65_2_groupi_n_24 & csa_tree_add_65_2_groupi_n_2)
    | ((csa_tree_add_65_2_groupi_n_2 & csa_tree_add_65_2_groupi_n_11) | (csa_tree_add_65_2_groupi_n_11 &
    csa_tree_add_65_2_groupi_n_24)));
 assign n_157 = (csa_tree_add_65_2_groupi_n_2 ^ (csa_tree_add_65_2_groupi_n_11 ^ csa_tree_add_65_2_groupi_n_24));
 assign csa_tree_add_65_2_groupi_n_24 = ((csa_tree_add_65_2_groupi_n_22 & csa_tree_add_65_2_groupi_n_12)
    | ((csa_tree_add_65_2_groupi_n_12 & csa_tree_add_65_2_groupi_n_3) | (csa_tree_add_65_2_groupi_n_3 & csa_tree_add_65_2_groupi_n_22)));
 assign n_158 = (csa_tree_add_65_2_groupi_n_12 ^ (csa_tree_add_65_2_groupi_n_3 ^ csa_tree_add_65_2_groupi_n_22));
 assign csa_tree_add_65_2_groupi_n_22 = ((csa_tree_add_65_2_groupi_n_20 & csa_tree_add_65_2_groupi_n_8)
    | ((csa_tree_add_65_2_groupi_n_8 & csa_tree_add_65_2_groupi_n_13) | (csa_tree_add_65_2_groupi_n_13 &
    csa_tree_add_65_2_groupi_n_20)));
 assign n_159 = (csa_tree_add_65_2_groupi_n_8 ^ (csa_tree_add_65_2_groupi_n_13 ^ csa_tree_add_65_2_groupi_n_20));
 assign csa_tree_add_65_2_groupi_n_20 = ((csa_tree_add_65_2_groupi_n_18 & csa_tree_add_65_2_groupi_n_6)
    | ((csa_tree_add_65_2_groupi_n_6 & csa_tree_add_65_2_groupi_n_9) | (csa_tree_add_65_2_groupi_n_9 & csa_tree_add_65_2_groupi_n_18)));
 assign n_160 = (csa_tree_add_65_2_groupi_n_6 ^ (csa_tree_add_65_2_groupi_n_9 ^ csa_tree_add_65_2_groupi_n_18));
 assign csa_tree_add_65_2_groupi_n_18 = ((csa_tree_add_65_2_groupi_n_16 & csa_tree_add_65_2_groupi_n_0)
    | ((csa_tree_add_65_2_groupi_n_0 & csa_tree_add_65_2_groupi_n_7) | (csa_tree_add_65_2_groupi_n_7 & csa_tree_add_65_2_groupi_n_16)));
 assign n_161 = (csa_tree_add_65_2_groupi_n_0 ^ (csa_tree_add_65_2_groupi_n_7 ^ csa_tree_add_65_2_groupi_n_16));
 assign csa_tree_add_65_2_groupi_n_16 = ((csa_tree_add_65_2_groupi_n_4 & {in8[1]}) | (({in8[1]} & csa_tree_add_65_2_groupi_n_1)
    | (csa_tree_add_65_2_groupi_n_1 & csa_tree_add_65_2_groupi_n_4)));
 assign n_162 = ({in8[1]} ^ (csa_tree_add_65_2_groupi_n_1 ^ csa_tree_add_65_2_groupi_n_4));
 assign csa_tree_add_65_2_groupi_n_14 = (({in7[7]} & {in6[7]}) | (({in6[7]} & {in8[7]}) | ({in8[7]} &
    {in7[7]})));
 assign csa_tree_add_65_2_groupi_n_15 = ({in6[7]} ^ ({in8[7]} ^ {in7[7]}));
 assign csa_tree_add_65_2_groupi_n_12 = (({in7[4]} & {in6[4]}) | (({in6[4]} & {in8[4]}) | ({in8[4]} &
    {in7[4]})));
 assign csa_tree_add_65_2_groupi_n_13 = ({in6[4]} ^ ({in8[4]} ^ {in7[4]}));
 assign csa_tree_add_65_2_groupi_n_10 = (({in7[6]} & {in6[6]}) | (({in6[6]} & {in8[6]}) | ({in8[6]} &
    {in7[6]})));
 assign csa_tree_add_65_2_groupi_n_11 = ({in6[6]} ^ ({in8[6]} ^ {in7[6]}));
 assign csa_tree_add_65_2_groupi_n_8 = (({in7[3]} & {in6[3]}) | (({in6[3]} & {in8[3]}) | ({in8[3]} &
    {in7[3]})));
 assign csa_tree_add_65_2_groupi_n_9 = ({in6[3]} ^ ({in8[3]} ^ {in7[3]}));
 assign csa_tree_add_65_2_groupi_n_6 = (({in7[2]} & {in6[2]}) | (({in6[2]} & {in8[2]}) | ({in8[2]} &
    {in7[2]})));
 assign csa_tree_add_65_2_groupi_n_7 = ({in6[2]} ^ ({in8[2]} ^ {in7[2]}));
 assign csa_tree_add_65_2_groupi_n_4 = (({in6[0]} & {in8[0]}) | (({in8[0]} & {in7[0]}) | ({in7[0]} &
    {in6[0]})));
 assign n_163 = ({in8[0]} ^ ({in7[0]} ^ {in6[0]}));
 assign csa_tree_add_65_2_groupi_n_2 = (({in8[5]} & {in6[5]}) | (({in6[5]} & {in7[5]}) | ({in7[5]} &
    {in8[5]})));
 assign csa_tree_add_65_2_groupi_n_3 = ({in6[5]} ^ ({in7[5]} ^ {in8[5]}));
 assign csa_tree_add_65_2_groupi_n_0 = ({in7[1]} & {in6[1]});
 assign csa_tree_add_65_2_groupi_n_1 = ({in7[1]} ^ {in6[1]});
 assign mul_71_11_n_263 = ((mul_71_11_n_184 & mul_71_11_n_209) | ((mul_71_11_n_209 & n_56) | (n_56 &
    mul_71_11_n_184)));
 assign mul_71_11_n_264 = (mul_71_11_n_209 ^ (n_56 ^ mul_71_11_n_184));
 assign mul_71_11_n_74 = ~((n_164 | mul_71_11_n_6) & (mul_71_11_n_27 | n_71));
 assign mul_71_11_n_99 = ~((n_164 | mul_71_11_n_7) & (mul_71_11_n_27 | n_61));
 assign mul_71_11_n_137 = ~(n_75 | mul_71_11_n_6);
 assign mul_71_11_n_43 = ~((n_164 | n_59) & (mul_71_11_n_27 | mul_71_11_n_20));
 assign mul_71_11_n_50 = ~((n_59 | n_74) & (mul_71_11_n_20 | mul_71_11_n_25));
 assign mul_71_11_n_101 = ~((n_71 | n_74) & (mul_71_11_n_6 | mul_71_11_n_25));
 assign mul_71_11_n_41 = ~((n_61 | n_74) & (mul_71_11_n_7 | mul_71_11_n_25));
 assign mul_71_11_n_102 = ~((n_56 | n_74) & (mul_71_11_n_19 | mul_71_11_n_25));
 assign mul_71_11_n_116 = ~((n_164 | n_56) & (mul_71_11_n_27 | mul_71_11_n_19));
 assign n_75 = ~(n_76 | (n_77 & mul_71_11_n_22));
 assign n_74 = ~mul_71_11_n_25;
 assign mul_71_11_n_278 = ((mul_71_11_n_174 & mul_71_11_n_215) | ((mul_71_11_n_215 & n_56) | (n_56 &
    mul_71_11_n_174)));
 assign mul_71_11_n_279 = (mul_71_11_n_215 ^ (n_56 ^ mul_71_11_n_174));
 assign mul_71_11_n_89 = ~((n_165 | n_71) & (mul_71_11_n_13 | mul_71_11_n_6));
 assign mul_71_11_n_83 = ~(n_77 & ~n_76);
 assign mul_71_11_n_186 = ~((mul_71_11_n_85 & n_165) | (mul_71_11_n_134 & n_60));
 assign mul_71_11_n_92 = ~((n_165 | n_61) & (mul_71_11_n_13 | mul_71_11_n_7));
 assign mul_71_11_n_79 = ~((n_71 & ~n_69) | (mul_71_11_n_6 & n_69));
 assign n_164 = ~(n_79 ^ n_68);
 assign mul_71_11_n_252 = ~((mul_71_11_n_121 & n_78) | (mul_71_11_n_145 & mul_71_11_n_22));
 assign mul_71_11_n_87 = ~((n_61 | n_62) & (mul_71_11_n_7 | mul_71_11_n_12));
 assign mul_71_11_n_67 = ~((n_71 | n_62) & (mul_71_11_n_6 | mul_71_11_n_12));
 assign mul_71_11_n_45 = ~((n_59 | n_62) & (mul_71_11_n_20 | mul_71_11_n_12));
 assign mul_71_11_n_112 = ~((n_56 | n_62) & (mul_71_11_n_19 | mul_71_11_n_12));
 assign mul_71_11_n_123 = ~((n_165 | n_56) & (mul_71_11_n_13 | mul_71_11_n_19));
 assign mul_71_11_n_42 = ~((n_165 | n_59) & (mul_71_11_n_13 | mul_71_11_n_20));
 assign n_76 = ~(n_69 | n_56);
 assign mul_71_11_n_251 = ~((mul_71_11_n_113 & mul_71_11_n_145) | (mul_71_11_n_103 & n_78));
 assign n_77 = ~(n_56 & n_69);
 assign mul_71_11_n_12 = ~n_62;
 assign n_79 = ((n_66 & n_67) | ((n_67 & n_58) | (n_58 & n_66)));
 assign n_165 = (n_67 ^ (n_58 ^ n_66));
 assign mul_71_11_n_118 = ~((n_56 | n_7) & (mul_71_11_n_19 | mul_71_11_n_16));
 assign mul_71_11_n_111 = ~((n_56 | n_16) & (mul_71_11_n_19 | mul_71_11_n_29));
 assign mul_71_11_n_104 = ~((n_56 | n_17) & (mul_71_11_n_19 | mul_71_11_n_28));
 assign mul_71_11_n_119 = ~((n_56 | n_6) & (mul_71_11_n_19 | mul_71_11_n_10));
 assign mul_71_11_n_114 = ~((n_56 | n_5) & (mul_71_11_n_19 | mul_71_11_n_26));
 assign mul_71_11_n_115 = ~((n_56 | n_14) & (mul_71_11_n_19 | mul_71_11_n_24));
 assign mul_71_11_n_117 = ~((n_56 | n_72) & (mul_71_11_n_19 | mul_71_11_n_15));
 assign mul_71_11_n_107 = ~((n_56 | n_18) & (mul_71_11_n_19 | mul_71_11_n_17));
 assign mul_71_11_n_120 = ~((n_56 | n_8) & (mul_71_11_n_19 | mul_71_11_n_14));
 assign mul_71_11_n_105 = ~((n_56 | n_11) & (mul_71_11_n_19 | mul_71_11_n_8));
 assign mul_71_11_n_109 = ~((n_56 | n_63) & (mul_71_11_n_19 | mul_71_11_n_30));
 assign mul_71_11_n_108 = ~((n_56 | n_73) & (mul_71_11_n_19 | mul_71_11_n_9));
 assign mul_71_11_n_106 = ~((n_56 | n_60) & (mul_71_11_n_19 | mul_71_11_n_11));
 assign mul_71_11_n_110 = ~((n_56 | n_12) & (mul_71_11_n_19 | mul_71_11_n_18));
 assign mul_71_11_n_121 = ~((n_56 | mul_71_11_n_23) & (mul_71_11_n_19 | n_64));
 assign n_0 = ~mul_68_11_n_246;
 assign mul_68_11_n_246 = ((n_167 & mul_68_11_n_155) | ((mul_68_11_n_155 & mul_68_11_n_185) | (mul_68_11_n_185
    & n_167)));
 assign n_2 = (mul_68_11_n_155 ^ (mul_68_11_n_185 ^ n_167));
 assign mul_71_11_n_145 = ~(n_78 | mul_71_11_n_19);
 assign n_1 = ~(add_51_2_n_15 ^ add_51_2_n_26);
 assign mul_71_11_n_19 = ~n_56;
 assign add_51_2_n_26 = (({in1[1]} & n_181) | ((n_181 & {in2[1]}) | ({in2[1]} & {in1[1]})));
 assign n_21 = (n_181 ^ ({in2[1]} ^ {in1[1]}));
 assign mul_71_11_n_124 = ~((n_61 | n_63) & (mul_71_11_n_7 | mul_71_11_n_30));
 assign mul_71_11_n_95 = ~((n_71 | n_63) & (mul_71_11_n_6 | mul_71_11_n_30));
 assign mul_71_11_n_57 = ~((n_59 | n_63) & (mul_71_11_n_20 | mul_71_11_n_30));
 assign mul_71_11_n_248 = ~(n_3 | mul_71_11_n_7);
 assign mul_71_11_n_247 = ~(n_4 | mul_71_11_n_20);
 assign n_13 = ~(n_23 ^ mul_68_11_n_189);
 assign mul_71_11_n_30 = ~n_63;
 assign n_3 = ~(n_9 | (n_10 & mul_71_11_n_22));
 assign n_4 = ~(n_19 | (n_20 & mul_71_11_n_22));
 assign mul_71_11_n_86 = ~(mul_71_11_n_135 & (n_59 | n_57));
 assign n_23 = ((mul_68_11_n_3 & mul_68_11_n_212) | ((mul_68_11_n_212 & mul_68_11_n_27) | (mul_68_11_n_27
    & mul_68_11_n_3)));
 assign n_22 = (mul_68_11_n_212 ^ (mul_68_11_n_27 ^ mul_68_11_n_3));
 assign n_24 = ((mul_68_11_n_200 & mul_68_11_n_213) | ((mul_68_11_n_213 & mul_68_11_n_104) | (mul_68_11_n_104
    & mul_68_11_n_200)));
 assign mul_68_11_n_266 = (mul_68_11_n_213 ^ (mul_68_11_n_104 ^ mul_68_11_n_200));
 assign n_167 = ((mul_68_11_n_176 & mul_68_11_n_178) | ((mul_68_11_n_178 & mul_68_11_n_116) | (mul_68_11_n_116
    & mul_68_11_n_176)));
 assign n_166 = (mul_68_11_n_178 ^ (mul_68_11_n_116 ^ mul_68_11_n_176));
 assign mul_71_11_n_81 = ~(n_20 & ~n_19);
 assign mul_71_11_n_84 = ~(n_10 & ~n_9);
 assign mul_71_11_n_237 = ~(mul_71_11_n_141 | (mul_71_11_n_143 & n_59));
 assign mul_71_11_n_185 = ~(mul_71_11_n_129 | (mul_71_11_n_130 & n_71));
 assign mul_71_11_n_241 = ~(mul_71_11_n_138 | (mul_71_11_n_139 & n_61));
 assign mul_71_11_n_56 = ~((n_59 | n_11) & (mul_71_11_n_20 | mul_71_11_n_8));
 assign mul_71_11_n_188 = ~((mul_71_11_n_85 & n_73) | (mul_71_11_n_134 & n_72));
 assign mul_71_11_n_78 = ~((n_59 & ~n_70) | (mul_71_11_n_20 & n_70));
 assign mul_71_11_n_80 = ~((n_61 & ~n_65) | (mul_71_11_n_7 & n_65));
 assign mul_71_11_n_127 = ~((n_61 | n_11) & (mul_71_11_n_7 | mul_71_11_n_8));
 assign mul_71_11_n_98 = ~((n_61 | n_5) & (mul_71_11_n_7 | mul_71_11_n_26));
 assign mul_71_11_n_97 = ~((n_61 | n_6) & (mul_71_11_n_7 | mul_71_11_n_10));
 assign mul_71_11_n_96 = ~((n_61 | n_14) & (mul_71_11_n_7 | mul_71_11_n_24));
 assign mul_71_11_n_72 = ~((n_61 | n_64) & (mul_71_11_n_7 | mul_71_11_n_23));
 assign mul_71_11_n_71 = ~((n_71 | n_14) & (mul_71_11_n_6 | mul_71_11_n_24));
 assign mul_71_11_n_70 = ~((n_61 | n_12) & (mul_71_11_n_7 | mul_71_11_n_18));
 assign mul_71_11_n_61 = ~((n_59 | n_14) & (mul_71_11_n_20 | mul_71_11_n_24));
 assign mul_71_11_n_38 = ~((n_61 | n_7) & (mul_71_11_n_7 | mul_71_11_n_16));
 assign mul_71_11_n_37 = ~((n_61 | n_8) & (mul_71_11_n_7 | mul_71_11_n_14));
 assign mul_71_11_n_88 = ~((n_71 | n_6) & (mul_71_11_n_6 | mul_71_11_n_10));
 assign mul_71_11_n_73 = ~((n_71 | n_7) & (mul_71_11_n_6 | mul_71_11_n_16));
 assign mul_71_11_n_60 = ~((n_59 | n_12) & (mul_71_11_n_20 | mul_71_11_n_18));
 assign mul_71_11_n_94 = ~((n_71 | n_64) & (mul_71_11_n_6 | mul_71_11_n_23));
 assign mul_71_11_n_59 = ~((n_59 | n_8) & (mul_71_11_n_20 | mul_71_11_n_14));
 assign mul_71_11_n_63 = ~((n_71 | n_8) & (mul_71_11_n_6 | mul_71_11_n_14));
 assign mul_71_11_n_40 = ~((n_71 | n_11) & (mul_71_11_n_6 | mul_71_11_n_8));
 assign mul_71_11_n_135 = ~(n_59 & n_57);
 assign mul_71_11_n_55 = ~((n_59 | n_16) & (mul_71_11_n_20 | mul_71_11_n_29));
 assign mul_71_11_n_54 = ~((n_59 | n_5) & (mul_71_11_n_20 | mul_71_11_n_26));
 assign mul_71_11_n_125 = ~((n_71 | n_5) & (mul_71_11_n_6 | mul_71_11_n_26));
 assign mul_71_11_n_53 = ~((n_59 | n_7) & (mul_71_11_n_20 | mul_71_11_n_16));
 assign mul_71_11_n_52 = ~((n_59 | n_18) & (mul_71_11_n_20 | mul_71_11_n_17));
 assign mul_71_11_n_39 = ~((n_71 | n_12) & (mul_71_11_n_6 | mul_71_11_n_18));
 assign mul_71_11_n_48 = ~((n_59 | n_64) & (mul_71_11_n_20 | mul_71_11_n_23));
 assign mul_71_11_n_47 = ~((n_59 | n_17) & (mul_71_11_n_20 | mul_71_11_n_28));
 assign mul_71_11_n_46 = ~((n_59 | n_6) & (mul_71_11_n_20 | mul_71_11_n_10));
 assign mul_71_11_n_100 = ~((n_61 | n_16) & (mul_71_11_n_7 | mul_71_11_n_29));
 assign mul_71_11_n_68 = ~((n_71 | n_16) & (mul_71_11_n_6 | mul_71_11_n_29));
 assign mul_71_11_n_69 = ~((n_61 | n_18) & (mul_71_11_n_7 | mul_71_11_n_17));
 assign mul_71_11_n_66 = ~((n_71 | n_18) & (mul_71_11_n_6 | mul_71_11_n_17));
 assign mul_71_11_n_126 = ~((n_71 | n_17) & (mul_71_11_n_6 | mul_71_11_n_28));
 assign mul_71_11_n_65 = ~((n_61 | n_17) & (mul_71_11_n_7 | mul_71_11_n_28));
 assign mul_71_11_n_91 = ~((n_61 | n_73) & (mul_71_11_n_7 | mul_71_11_n_9));
 assign mul_71_11_n_75 = ~((n_61 | n_72) & (mul_71_11_n_7 | mul_71_11_n_15));
 assign mul_71_11_n_58 = ~((n_59 | n_73) & (mul_71_11_n_20 | mul_71_11_n_9));
 assign mul_71_11_n_77 = ~((n_71 | n_72) & (mul_71_11_n_6 | mul_71_11_n_15));
 assign mul_71_11_n_76 = ~((n_71 | n_73) & (mul_71_11_n_6 | mul_71_11_n_9));
 assign mul_71_11_n_51 = ~((n_59 | n_72) & (mul_71_11_n_20 | mul_71_11_n_15));
 assign mul_71_11_n_49 = ~((n_59 | n_60) & (mul_71_11_n_20 | mul_71_11_n_11));
 assign mul_71_11_n_64 = ~((n_71 | n_60) & (mul_71_11_n_6 | mul_71_11_n_11));
 assign mul_71_11_n_62 = ~((n_61 | n_60) & (mul_71_11_n_7 | mul_71_11_n_11));
 assign mul_71_11_n_35 = ~((n_61 | n_15) & (mul_71_11_n_7 | mul_71_11_n_22));
 assign mul_71_11_n_33 = ~((n_59 | n_15) & (mul_71_11_n_20 | mul_71_11_n_22));
 assign mul_71_11_n_36 = ~((n_71 | n_15) & (mul_71_11_n_6 | mul_71_11_n_22));
 assign n_78 = ~mul_71_11_n_21;
 assign n_9 = ~(n_71 | n_65);
 assign n_10 = ~(n_65 & n_71);
 assign n_20 = ~(n_61 & n_70);
 assign n_19 = ~(n_70 | n_61);
 assign n_7 = ~mul_71_11_n_16;
 assign mul_71_11_n_23 = ~n_64;
 assign n_6 = ~mul_71_11_n_10;
 assign n_17 = ~mul_71_11_n_28;
 assign n_5 = ~mul_71_11_n_26;
 assign mul_71_11_n_9 = ~n_73;
 assign mul_71_11_n_7 = ~n_61;
 assign mul_71_11_n_20 = ~n_59;
 assign n_16 = ~mul_71_11_n_29;
 assign n_8 = ~mul_71_11_n_14;
 assign n_11 = ~mul_71_11_n_8;
 assign n_14 = ~mul_71_11_n_24;
 assign n_12 = ~mul_71_11_n_18;
 assign n_18 = ~mul_71_11_n_17;
 assign mul_71_11_n_11 = ~n_60;
 assign mul_71_11_n_15 = ~n_72;
 assign mul_71_11_n_6 = ~n_71;
 assign n_168 = ~(add_51_2_n_36 & (add_51_2_n_24 & (add_51_2_n_8 | add_51_2_n_6)));
 assign n_15 = ~mul_71_11_n_22;
 assign n_169 = ~(add_51_2_n_31 ^ add_51_2_n_20);
 assign n_170 = ~(mul_68_11_n_276 & (mul_68_11_n_358 | mul_68_11_n_279));
 assign n_171 = ~(mul_68_11_n_178 | (mul_68_11_n_177 & mul_68_11_n_94));
 assign n_172 = ~(add_51_2_n_28 ^ add_51_2_n_19);
 assign n_173 = ~(add_51_2_n_34 ^ add_51_2_n_14);
 assign n_174 = ~(mul_68_11_n_352 ^ mul_68_11_n_302);
 assign n_180 = ~(add_51_2_n_35 ^ add_51_2_n_13);
 assign n_175 = ~(mul_68_11_n_355 ^ mul_68_11_n_334);
 assign n_179 = ~(add_51_2_n_40 ^ add_51_2_n_17);
 assign n_176 = ~(mul_68_11_n_357 ^ mul_68_11_n_285);
 assign n_178 = ~({in2[0]} ^ {in1[0]});
 assign n_182 = ~n_177;
 assign n_177 = ~(n_153 & n_163);
 assign n_181 = ({in2[0]} & {in1[0]});
 assign n_184 = ~mul_68_11_n_351;
 assign n_187 = ~mul_68_11_n_283;
 assign n_25 = ~mul_68_11_n_255;
 assign n_186 = ~mul_68_11_n_290;
 assign n_183 = ~mul_68_11_n_332;
 assign n_188 = ~mul_68_11_n_331;
 assign n_189 = ~mul_68_11_n_311;
 assign n_185 = ~mul_68_11_n_319;
 assign n_190 = ~mul_68_11_n_273;
 assign n_191 = ~mul_68_11_n_292;
 assign mul_68_11_n_3 = (mul_68_11_n_105 | (mul_68_11_n_107 & mul_68_11_n_75));
 assign mul_68_11_n_358 = (mul_68_11_n_296 & (mul_68_11_n_352 | mul_68_11_n_297));
 assign mul_68_11_n_357 = ~(mul_68_11_n_296 & (mul_68_11_n_352 | mul_68_11_n_297));
 assign mul_68_11_n_355 = ~(mul_68_11_n_325 & (mul_68_11_n_351 | mul_68_11_n_327));
 assign mul_68_11_n_352 = ~(mul_68_11_n_349 | ~(mul_68_11_n_343 | mul_68_11_n_342));
 assign mul_68_11_n_351 = ~(mul_68_11_n_341 | (mul_68_11_n_347 & mul_68_11_n_337));
 assign mul_68_11_n_350 = ~(mul_68_11_n_321 & ~(mul_68_11_n_347 & mul_68_11_n_324));
 assign mul_68_11_n_349 = ~(mul_68_11_n_329 & (mul_68_11_n_346 & (mul_68_11_n_344 | mul_68_11_n_343)));
 assign mul_68_11_n_347 = ~(mul_68_11_n_344 & mul_68_11_n_342);
 assign mul_68_11_n_346 = ~(mul_68_11_n_330 | (mul_68_11_n_341 & mul_68_11_n_335));
 assign mul_68_11_n_344 = ~(mul_68_11_n_328 | ((mul_68_11_n_336 & mul_68_11_n_295) | (mul_68_11_n_326
    & mul_68_11_n_305)));
 assign mul_68_11_n_343 = ~(mul_68_11_n_337 & mul_68_11_n_335);
 assign mul_68_11_n_342 = ~(mul_68_11_n_310 & mul_68_11_n_336);
 assign mul_68_11_n_341 = ~(mul_68_11_n_312 & (mul_68_11_n_313 | mul_68_11_n_321));
 assign mul_68_11_n_340 = ~(mul_68_11_n_304 & (mul_68_11_n_322 | mul_68_11_n_303));
 assign mul_68_11_n_337 = ~(mul_68_11_n_313 | ~mul_68_11_n_324);
 assign mul_68_11_n_336 = ~(mul_68_11_n_303 | ~mul_68_11_n_326);
 assign mul_68_11_n_335 = ~(mul_68_11_n_327 | mul_68_11_n_323);
 assign mul_68_11_n_334 = ~(mul_68_11_n_329 & ~mul_68_11_n_323);
 assign mul_68_11_n_333 = ~(mul_68_11_n_327 | ~mul_68_11_n_325);
 assign mul_68_11_n_332 = ~(mul_68_11_n_324 & mul_68_11_n_321);
 assign mul_68_11_n_331 = ~(mul_68_11_n_326 & ~mul_68_11_n_328);
 assign mul_68_11_n_330 = ~(mul_68_11_n_325 | mul_68_11_n_323);
 assign mul_68_11_n_329 = ~(mul_68_11_n_294 & mul_68_11_n_316);
 assign mul_68_11_n_328 = (mul_68_11_n_315 & mul_68_11_n_298);
 assign mul_68_11_n_327 = ~(mul_68_11_n_317 | mul_68_11_n_308);
 assign mul_68_11_n_326 = (mul_68_11_n_315 | mul_68_11_n_298);
 assign mul_68_11_n_325 = ~(mul_68_11_n_317 & mul_68_11_n_308);
 assign mul_68_11_n_324 = (mul_68_11_n_307 | mul_68_11_n_314);
 assign mul_68_11_n_319 = ~(mul_68_11_n_312 & ~mul_68_11_n_313);
 assign mul_68_11_n_318 = ~(mul_68_11_n_278 & (mul_68_11_n_301 | mul_68_11_n_277));
 assign mul_68_11_n_323 = ~(mul_68_11_n_294 | mul_68_11_n_316);
 assign mul_68_11_n_322 = ~(mul_68_11_n_310 | mul_68_11_n_295);
 assign mul_68_11_n_321 = ~(mul_68_11_n_307 & mul_68_11_n_314);
 assign mul_68_11_n_316 = ((mul_68_11_n_258 & mul_68_11_n_264) | ((mul_68_11_n_264 & mul_68_11_n_227)
    | (mul_68_11_n_227 & mul_68_11_n_258)));
 assign mul_68_11_n_317 = (mul_68_11_n_264 ^ (mul_68_11_n_227 ^ mul_68_11_n_258));
 assign mul_68_11_n_314 = ((mul_68_11_n_252 & mul_68_11_n_225) | ((mul_68_11_n_225 & mul_68_11_n_260)
    | (mul_68_11_n_260 & mul_68_11_n_252)));
 assign mul_68_11_n_315 = (mul_68_11_n_225 ^ (mul_68_11_n_260 ^ mul_68_11_n_252));
 assign mul_68_11_n_313 = ~(mul_68_11_n_309 | mul_68_11_n_306);
 assign mul_68_11_n_312 = ~(mul_68_11_n_309 & mul_68_11_n_306);
 assign mul_68_11_n_311 = ~(mul_68_11_n_303 | mul_68_11_n_305);
 assign mul_68_11_n_310 = ~(mul_68_11_n_287 | (mul_68_11_n_277 | mul_68_11_n_301));
 assign mul_68_11_n_308 = ((mul_68_11_n_259 & mul_68_11_n_203) | ((mul_68_11_n_203 & mul_68_11_n_253)
    | (mul_68_11_n_253 & mul_68_11_n_259)));
 assign mul_68_11_n_309 = (mul_68_11_n_203 ^ (mul_68_11_n_253 ^ mul_68_11_n_259));
 assign mul_68_11_n_306 = ((mul_68_11_n_251 & mul_68_11_n_254) | ((mul_68_11_n_254 & mul_68_11_n_195)
    | (mul_68_11_n_195 & mul_68_11_n_251)));
 assign mul_68_11_n_307 = (mul_68_11_n_254 ^ (mul_68_11_n_195 ^ mul_68_11_n_251));
 assign mul_68_11_n_305 = ~mul_68_11_n_304;
 assign mul_68_11_n_304 = ~(mul_68_11_n_299 & mul_68_11_n_280);
 assign mul_68_11_n_303 = ~(mul_68_11_n_299 | mul_68_11_n_280);
 assign mul_68_11_n_302 = ~(mul_68_11_n_297 | ~mul_68_11_n_296);
 assign mul_68_11_n_301 = ~(mul_68_11_n_291 | ((mul_68_11_n_286 & mul_68_11_n_265) | (mul_68_11_n_286
    & mul_68_11_n_240)));
 assign mul_68_11_n_298 = ((mul_68_11_n_261 & mul_68_11_n_205) | ((mul_68_11_n_205 & mul_68_11_n_241)
    | (mul_68_11_n_241 & mul_68_11_n_261)));
 assign mul_68_11_n_299 = (mul_68_11_n_205 ^ (mul_68_11_n_241 ^ mul_68_11_n_261));
 assign mul_68_11_n_297 = ~(mul_68_11_n_268 | mul_68_11_n_293);
 assign mul_68_11_n_296 = ~(mul_68_11_n_268 & mul_68_11_n_293);
 assign mul_68_11_n_295 = ~(mul_68_11_n_288 & (mul_68_11_n_287 | mul_68_11_n_278));
 assign mul_68_11_n_293 = ((mul_68_11_n_263 & mul_68_11_n_226) | ((mul_68_11_n_226 & mul_68_11_n_235)
    | (mul_68_11_n_235 & mul_68_11_n_263)));
 assign mul_68_11_n_294 = (mul_68_11_n_226 ^ (mul_68_11_n_235 ^ mul_68_11_n_263));
 assign mul_68_11_n_292 = ~(mul_68_11_n_288 & ~mul_68_11_n_287);
 assign mul_68_11_n_291 = ~(mul_68_11_n_274 & (mul_68_11_n_275 | mul_68_11_n_248));
 assign mul_68_11_n_290 = ~(mul_68_11_n_248 & (mul_68_11_n_273 | mul_68_11_n_249));
 assign mul_68_11_n_288 = ~(mul_68_11_n_281 & mul_68_11_n_271);
 assign mul_68_11_n_287 = ~(mul_68_11_n_281 | mul_68_11_n_271);
 assign mul_68_11_n_286 = ~(mul_68_11_n_275 | mul_68_11_n_249);
 assign mul_68_11_n_285 = ~(mul_68_11_n_276 & ~mul_68_11_n_279);
 assign mul_68_11_n_284 = ~(mul_68_11_n_274 & ~mul_68_11_n_275);
 assign mul_68_11_n_283 = ~(mul_68_11_n_277 | ~mul_68_11_n_278);
 assign mul_68_11_n_280 = ((mul_68_11_n_242 & mul_68_11_n_214) | ((mul_68_11_n_214 & mul_68_11_n_199)
    | (mul_68_11_n_199 & mul_68_11_n_242)));
 assign mul_68_11_n_281 = (mul_68_11_n_214 ^ (mul_68_11_n_199 ^ mul_68_11_n_242));
 assign mul_68_11_n_279 = ~(mul_68_11_n_266 | mul_68_11_n_267);
 assign mul_68_11_n_278 = ~(mul_68_11_n_272 & mul_68_11_n_269);
 assign mul_68_11_n_277 = ~(mul_68_11_n_272 | mul_68_11_n_269);
 assign mul_68_11_n_276 = ~(mul_68_11_n_266 & mul_68_11_n_267);
 assign mul_68_11_n_275 = ~(mul_68_11_n_270 | mul_68_11_n_243);
 assign mul_68_11_n_274 = ~(mul_68_11_n_270 & mul_68_11_n_243);
 assign mul_68_11_n_273 = ~(mul_68_11_n_240 | mul_68_11_n_265);
 assign mul_68_11_n_271 = ((mul_68_11_n_222 & mul_68_11_n_215) | ((mul_68_11_n_215 & mul_68_11_n_217)
    | (mul_68_11_n_217 & mul_68_11_n_222)));
 assign mul_68_11_n_272 = (mul_68_11_n_215 ^ (mul_68_11_n_217 ^ mul_68_11_n_222));
 assign mul_68_11_n_263 = ((mul_68_11_n_202 & mul_68_11_n_208) | ((mul_68_11_n_208 & mul_68_11_n_26)
    | (mul_68_11_n_26 & mul_68_11_n_202)));
 assign mul_68_11_n_264 = (mul_68_11_n_208 ^ (mul_68_11_n_26 ^ mul_68_11_n_202));
 assign mul_68_11_n_269 = ((mul_68_11_n_223 & mul_68_11_n_187) | ((mul_68_11_n_187 & mul_68_11_n_210)
    | (mul_68_11_n_210 & mul_68_11_n_223)));
 assign mul_68_11_n_270 = (mul_68_11_n_187 ^ (mul_68_11_n_210 ^ mul_68_11_n_223));
 assign mul_68_11_n_267 = ((mul_68_11_n_234 & mul_68_11_n_190) | ((mul_68_11_n_190 & mul_68_11_n_201)
    | (mul_68_11_n_201 & mul_68_11_n_234)));
 assign mul_68_11_n_268 = (mul_68_11_n_190 ^ (mul_68_11_n_201 ^ mul_68_11_n_234));
 assign mul_68_11_n_260 = ((mul_68_11_n_198 & mul_68_11_n_207) | ((mul_68_11_n_207 & mul_68_11_n_181)
    | (mul_68_11_n_181 & mul_68_11_n_198)));
 assign mul_68_11_n_261 = (mul_68_11_n_207 ^ (mul_68_11_n_181 ^ mul_68_11_n_198));
 assign mul_68_11_n_258 = ((mul_68_11_n_194 & mul_68_11_n_196) | ((mul_68_11_n_196 & mul_68_11_n_209)
    | (mul_68_11_n_209 & mul_68_11_n_194)));
 assign mul_68_11_n_259 = (mul_68_11_n_196 ^ (mul_68_11_n_209 ^ mul_68_11_n_194));
 assign mul_68_11_n_265 = ~(mul_68_11_n_250 | mul_68_11_n_233);
 assign mul_68_11_n_257 = ~(mul_68_11_n_249 | ~mul_68_11_n_248);
 assign mul_68_11_n_255 = ~(mul_68_11_n_250 & mul_68_11_n_230);
 assign mul_68_11_n_253 = ((mul_68_11_n_197 & mul_68_11_n_224) | ((mul_68_11_n_224 & mul_68_11_n_192)
    | (mul_68_11_n_192 & mul_68_11_n_197)));
 assign mul_68_11_n_254 = (mul_68_11_n_224 ^ (mul_68_11_n_192 ^ mul_68_11_n_197));
 assign mul_68_11_n_251 = ((mul_68_11_n_193 & mul_68_11_n_206) | ((mul_68_11_n_206 & mul_68_11_n_204)
    | (mul_68_11_n_204 & mul_68_11_n_193)));
 assign mul_68_11_n_252 = (mul_68_11_n_206 ^ (mul_68_11_n_204 ^ mul_68_11_n_193));
 assign mul_68_11_n_250 = ~(mul_68_11_n_246 & ~mul_68_11_n_232);
 assign mul_68_11_n_249 = ~(mul_68_11_n_244 | mul_68_11_n_220);
 assign mul_68_11_n_248 = ~(mul_68_11_n_244 & mul_68_11_n_220);
 assign mul_68_11_n_243 = ((mul_68_11_n_211 & mul_68_11_n_183) | ((mul_68_11_n_183 & mul_68_11_n_123)
    | (mul_68_11_n_123 & mul_68_11_n_211)));
 assign mul_68_11_n_244 = (mul_68_11_n_183 ^ (mul_68_11_n_123 ^ mul_68_11_n_211));
 assign mul_68_11_n_241 = ((mul_68_11_n_216 & mul_68_11_n_182) | ((mul_68_11_n_182 & mul_68_11_n_157)
    | (mul_68_11_n_157 & mul_68_11_n_216)));
 assign mul_68_11_n_242 = (mul_68_11_n_182 ^ (mul_68_11_n_157 ^ mul_68_11_n_216));
 assign mul_68_11_n_240 = ~(mul_68_11_n_231 & (mul_68_11_n_233 | mul_68_11_n_230));
 assign mul_68_11_n_237 = ~(mul_68_11_n_231 & ~mul_68_11_n_233);
 assign mul_68_11_n_236 = ~(mul_68_11_n_230 & ~mul_68_11_n_232);
 assign mul_68_11_n_234 = ((mul_68_11_n_191 & mul_68_11_n_103) | ((mul_68_11_n_103 & mul_68_11_n_158)
    | (mul_68_11_n_158 & mul_68_11_n_191)));
 assign mul_68_11_n_235 = (mul_68_11_n_103 ^ (mul_68_11_n_158 ^ mul_68_11_n_191));
 assign mul_68_11_n_233 = ~(mul_68_11_n_221 | mul_68_11_n_228);
 assign mul_68_11_n_232 = ~(mul_68_11_n_229 | mul_68_11_n_188);
 assign mul_68_11_n_231 = ~(mul_68_11_n_221 & mul_68_11_n_228);
 assign mul_68_11_n_230 = ~(mul_68_11_n_229 & mul_68_11_n_188);
 assign mul_68_11_n_228 = ((mul_68_11_n_151 & mul_68_11_n_162) | ((mul_68_11_n_162 & mul_68_11_n_100)
    | (mul_68_11_n_100 & mul_68_11_n_151)));
 assign mul_68_11_n_229 = (mul_68_11_n_162 ^ (mul_68_11_n_100 ^ mul_68_11_n_151));
 assign mul_68_11_n_226 = ((mul_68_11_n_147 & mul_68_11_n_128) | ((mul_68_11_n_128 & mul_68_11_n_139)
    | (mul_68_11_n_139 & mul_68_11_n_147)));
 assign mul_68_11_n_227 = (mul_68_11_n_128 ^ (mul_68_11_n_139 ^ mul_68_11_n_147));
 assign mul_68_11_n_224 = ((mul_68_11_n_153 & mul_68_11_n_137) | ((mul_68_11_n_137 & mul_68_11_n_138)
    | (mul_68_11_n_138 & mul_68_11_n_153)));
 assign mul_68_11_n_225 = (mul_68_11_n_137 ^ (mul_68_11_n_138 ^ mul_68_11_n_153));
 assign mul_68_11_n_222 = ((mul_68_11_n_154 & mul_68_11_n_156) | ((mul_68_11_n_156 & mul_68_11_n_127)
    | (mul_68_11_n_127 & mul_68_11_n_154)));
 assign mul_68_11_n_223 = (mul_68_11_n_156 ^ (mul_68_11_n_127 ^ mul_68_11_n_154));
 assign mul_68_11_n_220 = ((mul_68_11_n_184 & mul_68_11_n_124) | ((mul_68_11_n_124 & mul_68_11_n_161)
    | (mul_68_11_n_161 & mul_68_11_n_184)));
 assign mul_68_11_n_221 = (mul_68_11_n_124 ^ (mul_68_11_n_161 ^ mul_68_11_n_184));
 assign mul_68_11_n_216 = ((mul_68_11_n_130 & mul_68_11_n_118) | ((mul_68_11_n_118 & mul_68_11_n_164)
    | (mul_68_11_n_164 & mul_68_11_n_130)));
 assign mul_68_11_n_217 = (mul_68_11_n_118 ^ (mul_68_11_n_164 ^ mul_68_11_n_130));
 assign mul_68_11_n_214 = ((mul_68_11_n_186 & mul_68_11_n_142) | ((mul_68_11_n_142 & mul_68_11_n_160)
    | (mul_68_11_n_160 & mul_68_11_n_186)));
 assign mul_68_11_n_215 = (mul_68_11_n_142 ^ (mul_68_11_n_160 ^ mul_68_11_n_186));
 assign mul_68_11_n_212 = ((mul_68_11_n_144 & mul_68_11_n_22) | ((mul_68_11_n_22 & mul_68_11_n_159) |
    (mul_68_11_n_159 & mul_68_11_n_144)));
 assign mul_68_11_n_213 = (mul_68_11_n_22 ^ (mul_68_11_n_159 ^ mul_68_11_n_144));
 assign mul_68_11_n_210 = ((mul_68_11_n_152 & mul_68_11_n_165) | ((mul_68_11_n_165 & mul_68_11_n_117)
    | (mul_68_11_n_117 & mul_68_11_n_152)));
 assign mul_68_11_n_211 = (mul_68_11_n_165 ^ (mul_68_11_n_117 ^ mul_68_11_n_152));
 assign mul_68_11_n_208 = ((mul_68_11_n_174 & mul_68_11_n_121) | ((mul_68_11_n_121 & mul_68_11_n_11)
    | (mul_68_11_n_11 & mul_68_11_n_174)));
 assign mul_68_11_n_209 = (mul_68_11_n_121 ^ (mul_68_11_n_11 ^ mul_68_11_n_174));
 assign mul_68_11_n_206 = ((mul_68_11_n_166 & mul_68_11_n_122) | ((mul_68_11_n_122 & mul_68_11_n_21)
    | (mul_68_11_n_21 & mul_68_11_n_166)));
 assign mul_68_11_n_207 = (mul_68_11_n_122 ^ (mul_68_11_n_21 ^ mul_68_11_n_166));
 assign mul_68_11_n_204 = ((mul_68_11_n_145 & mul_68_11_n_135) | ((mul_68_11_n_135 & mul_68_11_n_132)
    | (mul_68_11_n_132 & mul_68_11_n_145)));
 assign mul_68_11_n_205 = (mul_68_11_n_135 ^ (mul_68_11_n_132 ^ mul_68_11_n_145));
 assign mul_68_11_n_202 = ((mul_68_11_n_148 & mul_68_11_n_29) | ((mul_68_11_n_29 & mul_68_11_n_134) |
    (mul_68_11_n_134 & mul_68_11_n_148)));
 assign mul_68_11_n_203 = (mul_68_11_n_29 ^ (mul_68_11_n_134 ^ mul_68_11_n_148));
 assign mul_68_11_n_200 = ((mul_68_11_n_172 & mul_68_11_n_140) | ((mul_68_11_n_140 & mul_68_11_n_30)
    | (mul_68_11_n_30 & mul_68_11_n_172)));
 assign mul_68_11_n_201 = (mul_68_11_n_140 ^ (mul_68_11_n_30 ^ mul_68_11_n_172));
 assign mul_68_11_n_198 = ((mul_68_11_n_146 & mul_68_11_n_133) | ((mul_68_11_n_133 & mul_68_11_n_163)
    | (mul_68_11_n_163 & mul_68_11_n_146)));
 assign mul_68_11_n_199 = (mul_68_11_n_133 ^ (mul_68_11_n_163 ^ mul_68_11_n_146));
 assign mul_68_11_n_196 = ((mul_68_11_n_167 & mul_68_11_n_129) | ((mul_68_11_n_129 & n_162) | (n_162
    & mul_68_11_n_167)));
 assign mul_68_11_n_197 = (mul_68_11_n_129 ^ (n_162 ^ mul_68_11_n_167));
 assign mul_68_11_n_194 = ((mul_68_11_n_168 & mul_68_11_n_23) | ((mul_68_11_n_23 & mul_68_11_n_141) |
    (mul_68_11_n_141 & mul_68_11_n_168)));
 assign mul_68_11_n_195 = (mul_68_11_n_23 ^ (mul_68_11_n_141 ^ mul_68_11_n_168));
 assign mul_68_11_n_192 = ((mul_68_11_n_126 & mul_68_11_n_28) | ((mul_68_11_n_28 & n_162) | (n_162 &
    mul_68_11_n_126)));
 assign mul_68_11_n_193 = (mul_68_11_n_28 ^ (n_162 ^ mul_68_11_n_126));
 assign mul_68_11_n_190 = ((mul_68_11_n_131 & mul_68_11_n_136) | ((mul_68_11_n_136 & mul_68_11_n_20)
    | (mul_68_11_n_20 & mul_68_11_n_131)));
 assign mul_68_11_n_191 = (mul_68_11_n_136 ^ (mul_68_11_n_20 ^ mul_68_11_n_131));
 assign mul_68_11_n_189 = ~(mul_68_11_n_179 ^ mul_68_11_n_27);
 assign mul_68_11_n_186 = (mul_68_11_n_149 & mul_68_11_n_171);
 assign mul_68_11_n_187 = (mul_68_11_n_149 ^ mul_68_11_n_171);
 assign mul_68_11_n_188 = (mul_68_11_n_173 & mul_68_11_n_170);
 assign mul_68_11_n_185 = (mul_68_11_n_173 ^ mul_68_11_n_170);
 assign mul_68_11_n_183 = (mul_68_11_n_150 & mul_68_11_n_143);
 assign mul_68_11_n_184 = (mul_68_11_n_150 ^ mul_68_11_n_143);
 assign mul_68_11_n_181 = (mul_68_11_n_125 & mul_68_11_n_169);
 assign mul_68_11_n_182 = (mul_68_11_n_125 ^ mul_68_11_n_169);
 assign mul_68_11_n_179 = ~(mul_68_11_n_175 ^ mul_68_11_n_24);
 assign mul_68_11_n_178 = ~(mul_68_11_n_177 | mul_68_11_n_94);
 assign mul_68_11_n_177 = ~((mul_68_11_n_119 & mul_68_11_n_33) | (mul_68_11_n_87 & n_163));
 assign mul_68_11_n_176 = ~((mul_68_11_n_120 | mul_68_11_n_88) & (mul_68_11_n_83 | mul_68_11_n_13));
 assign mul_68_11_n_175 = ~(mul_68_11_n_105 | (mul_68_11_n_107 & n_154));
 assign mul_68_11_n_174 = ~(mul_68_11_n_110 | (mul_68_11_n_114 & n_160));
 assign mul_68_11_n_173 = ~((mul_68_11_n_120 | mul_68_11_n_83) & (mul_68_11_n_81 | mul_68_11_n_13));
 assign mul_68_11_n_172 = ~(mul_68_11_n_109 & ~(mul_68_11_n_112 & mul_68_11_n_58));
 assign mul_68_11_n_171 = ~(mul_68_11_n_12 | ((mul_68_11_n_1 & n_153) | (n_158 & n_157)));
 assign mul_68_11_n_170 = ~(mul_68_11_n_5 | ((mul_68_11_n_0 & n_153) | (n_162 & n_161)));
 assign mul_68_11_n_169 = ~(mul_68_11_n_4 | ((mul_68_11_n_2 & n_153) | (n_156 & n_155)));
 assign mul_68_11_n_168 = ~((mul_68_11_n_113 | mul_68_11_n_50) & (mul_68_11_n_70 | mul_68_11_n_56));
 assign mul_68_11_n_167 = ~(mul_68_11_n_111 & ~(mul_68_11_n_114 & mul_68_11_n_39));
 assign mul_68_11_n_166 = ~((mul_68_11_n_120 | mul_68_11_n_82) & (mul_68_11_n_13 | mul_68_11_n_11));
 assign mul_68_11_n_165 = ~((mul_68_11_n_120 | mul_68_11_n_85) & (mul_68_11_n_86 | mul_68_11_n_13));
 assign mul_68_11_n_164 = ~((mul_68_11_n_115 | mul_68_11_n_42) & (mul_68_11_n_71 | mul_68_11_n_93));
 assign mul_68_11_n_163 = ~((mul_68_11_n_120 | mul_68_11_n_80) & (mul_68_11_n_82 | mul_68_11_n_13));
 assign mul_68_11_n_162 = ~((mul_68_11_n_120 | mul_68_11_n_81) & (mul_68_11_n_84 | mul_68_11_n_13));
 assign mul_68_11_n_161 = ~((mul_68_11_n_120 | mul_68_11_n_84) & (mul_68_11_n_85 | mul_68_11_n_13));
 assign mul_68_11_n_160 = ~((mul_68_11_n_120 | mul_68_11_n_89) & (mul_68_11_n_80 | mul_68_11_n_13));
 assign mul_68_11_n_159 = ~(mul_68_11_n_108 | (mul_68_11_n_112 & n_156));
 assign mul_68_11_n_158 = ~((mul_68_11_n_113 | mul_68_11_n_43) & (mul_68_11_n_70 | mul_68_11_n_57));
 assign mul_68_11_n_157 = ~((mul_68_11_n_113 | mul_68_11_n_45) & (mul_68_11_n_70 | mul_68_11_n_46));
 assign mul_68_11_n_156 = ~((mul_68_11_n_120 | mul_68_11_n_86) & (mul_68_11_n_89 | mul_68_11_n_13));
 assign mul_68_11_n_155 = ~((mul_68_11_n_115 | mul_68_11_n_36) & (mul_68_11_n_71 | mul_68_11_n_41));
 assign mul_68_11_n_154 = ~((mul_68_11_n_113 | mul_68_11_n_37) & (mul_68_11_n_70 | mul_68_11_n_63));
 assign mul_68_11_n_153 = ~((mul_68_11_n_113 | mul_68_11_n_60) & (mul_68_11_n_70 | mul_68_11_n_50));
 assign mul_68_11_n_152 = ~((mul_68_11_n_115 | mul_68_11_n_95) & (mul_68_11_n_71 | mul_68_11_n_61));
 assign mul_68_11_n_151 = ~((mul_68_11_n_115 | mul_68_11_n_41) & (mul_68_11_n_71 | mul_68_11_n_55));
 assign mul_68_11_n_150 = ~((mul_68_11_n_115 | mul_68_11_n_55) & (mul_68_11_n_71 | mul_68_11_n_95));
 assign mul_68_11_n_149 = ~((mul_68_11_n_115 | mul_68_11_n_61) & (mul_68_11_n_71 | mul_68_11_n_42));
 assign mul_68_11_n_148 = ~((mul_68_11_n_113 | mul_68_11_n_56) & (mul_68_11_n_70 | mul_68_11_n_54));
 assign mul_68_11_n_147 = ~((mul_68_11_n_113 | mul_68_11_n_54) & (mul_68_11_n_70 | mul_68_11_n_43));
 assign mul_68_11_n_146 = ~((mul_68_11_n_115 | mul_68_11_n_93) & (mul_68_11_n_71 | mul_68_11_n_48));
 assign mul_68_11_n_145 = ~((mul_68_11_n_106 | mul_68_11_n_77) & (mul_68_11_n_69 | mul_68_11_n_78));
 assign mul_68_11_n_144 = ((mul_68_11_n_102 & mul_68_11_n_75) | (mul_68_11_n_107 & mul_68_11_n_101));
 assign mul_68_11_n_143 = ~(mul_68_11_n_6 | ((mul_68_11_n_25 & n_159) | (n_160 & n_153)));
 assign mul_68_11_n_142 = ~((mul_68_11_n_113 | mul_68_11_n_63) & (mul_68_11_n_70 | mul_68_11_n_45));
 assign mul_68_11_n_141 = ~((mul_68_11_n_106 | mul_68_11_n_76) & (mul_68_11_n_69 | mul_68_11_n_74));
 assign mul_68_11_n_140 = ~((mul_68_11_n_106 | mul_68_11_n_79) & (mul_68_11_n_69 | mul_68_11_n_73));
 assign mul_68_11_n_139 = ~((mul_68_11_n_106 | mul_68_11_n_90) & (mul_68_11_n_69 | mul_68_11_n_72));
 assign mul_68_11_n_138 = ~((mul_68_11_n_106 | mul_68_11_n_78) & (mul_68_11_n_69 | mul_68_11_n_76));
 assign mul_68_11_n_137 = ~((mul_68_11_n_115 | mul_68_11_n_49) & (mul_68_11_n_71 | mul_68_11_n_38));
 assign mul_68_11_n_136 = ~((mul_68_11_n_106 | mul_68_11_n_72) & (mul_68_11_n_69 | mul_68_11_n_79));
 assign mul_68_11_n_135 = ~((mul_68_11_n_115 | mul_68_11_n_48) & (mul_68_11_n_71 | mul_68_11_n_49));
 assign mul_68_11_n_134 = ~((mul_68_11_n_106 | mul_68_11_n_74) & (mul_68_11_n_69 | mul_68_11_n_90));
 assign mul_68_11_n_133 = ~((mul_68_11_n_106 | mul_68_11_n_34) & (mul_68_11_n_69 | mul_68_11_n_77));
 assign mul_68_11_n_132 = ~((mul_68_11_n_113 | mul_68_11_n_46) & (mul_68_11_n_70 | mul_68_11_n_60));
 assign mul_68_11_n_131 = ~(mul_68_11_n_98 | (mul_68_11_n_96 & n_158));
 assign mul_68_11_n_130 = ~((mul_68_11_n_97 | mul_68_11_n_44) & (mul_68_11_n_68 | mul_68_11_n_52));
 assign mul_68_11_n_129 = ~((mul_68_11_n_97 | mul_68_11_n_53) & (mul_68_11_n_68 | mul_68_11_n_47));
 assign mul_68_11_n_128 = ~(mul_68_11_n_99 & ~(mul_68_11_n_96 & mul_68_11_n_92));
 assign mul_68_11_n_127 = ~((mul_68_11_n_97 | mul_68_11_n_62) & (mul_68_11_n_68 | mul_68_11_n_44));
 assign mul_68_11_n_126 = ~((mul_68_11_n_97 | mul_68_11_n_59) & (mul_68_11_n_68 | mul_68_11_n_53));
 assign mul_68_11_n_125 = ~((mul_68_11_n_97 | mul_68_11_n_52) & (mul_68_11_n_68 | mul_68_11_n_40));
 assign mul_68_11_n_124 = ~((mul_68_11_n_97 | mul_68_11_n_35) & (mul_68_11_n_68 | mul_68_11_n_51));
 assign mul_68_11_n_123 = ~((mul_68_11_n_97 | mul_68_11_n_51) & (mul_68_11_n_68 | mul_68_11_n_62));
 assign mul_68_11_n_122 = ~((mul_68_11_n_97 | mul_68_11_n_40) & (mul_68_11_n_68 | mul_68_11_n_59));
 assign mul_68_11_n_121 = ~((mul_68_11_n_97 | mul_68_11_n_47) & (mul_68_11_n_68 | mul_68_11_n_91));
 assign mul_68_11_n_119 = ~mul_68_11_n_120;
 assign mul_68_11_n_120 = ~(mul_68_11_n_32 & mul_68_11_n_13);
 assign mul_68_11_n_118 = ~(mul_68_11_n_69 | mul_68_11_n_7);
 assign mul_68_11_n_117 = ~(mul_68_11_n_70 | mul_68_11_n_7);
 assign mul_68_11_n_116 = ~(mul_68_11_n_71 | mul_68_11_n_7);
 assign mul_68_11_n_114 = ~mul_68_11_n_115;
 assign mul_68_11_n_115 = ~(mul_68_11_n_71 & mul_68_11_n_67);
 assign mul_68_11_n_112 = ~mul_68_11_n_113;
 assign mul_68_11_n_113 = ~(mul_68_11_n_70 & mul_68_11_n_66);
 assign mul_68_11_n_111 = ~mul_68_11_n_110;
 assign mul_68_11_n_110 = ~(mul_68_11_n_71 | mul_68_11_n_5);
 assign mul_68_11_n_109 = ~mul_68_11_n_108;
 assign mul_68_11_n_108 = ~(mul_68_11_n_70 | mul_68_11_n_12);
 assign mul_68_11_n_107 = ~mul_68_11_n_106;
 assign mul_68_11_n_106 = ~(mul_68_11_n_69 & mul_68_11_n_65);
 assign mul_68_11_n_105 = ~(mul_68_11_n_69 | mul_68_11_n_4);
 assign mul_68_11_n_104 = ~mul_68_11_n_30;
 assign mul_68_11_n_103 = ~mul_68_11_n_26;
 assign mul_68_11_n_102 = ~mul_68_11_n_69;
 assign mul_68_11_n_101 = ~mul_68_11_n_73;
 assign mul_68_11_n_100 = ~(mul_68_11_n_68 | mul_68_11_n_7);
 assign mul_68_11_n_99 = ~mul_68_11_n_98;
 assign mul_68_11_n_96 = ~mul_68_11_n_97;
 assign mul_68_11_n_98 = ~(mul_68_11_n_68 | mul_68_11_n_6);
 assign mul_68_11_n_97 = ~(mul_68_11_n_68 & mul_68_11_n_64);
 assign mul_68_11_n_92 = ~mul_68_11_n_91;
 assign mul_68_11_n_88 = ~mul_68_11_n_87;
 assign mul_68_11_n_67 = ~((mul_68_11_n_5 & ~n_161) | (n_160 & n_161));
 assign mul_68_11_n_66 = ~((mul_68_11_n_12 & ~n_157) | (n_156 & n_157));
 assign mul_68_11_n_65 = ~((mul_68_11_n_4 & ~n_155) | (n_154 & n_155));
 assign mul_68_11_n_64 = ~((mul_68_11_n_6 & ~n_159) | (n_158 & n_159));
 assign mul_68_11_n_95 = ~((mul_68_11_n_5 & n_150) | (mul_68_11_n_18 & n_160));
 assign mul_68_11_n_94 = ~(n_162 & ~n_182);
 assign mul_68_11_n_93 = ~((mul_68_11_n_5 & n_147) | (mul_68_11_n_16 & n_160));
 assign mul_68_11_n_91 = ~((mul_68_11_n_6 & n_144) | (mul_68_11_n_15 & n_158));
 assign mul_68_11_n_90 = ~((mul_68_11_n_4 & n_148) | (mul_68_11_n_9 & n_154));
 assign mul_68_11_n_89 = ~((mul_68_11_n_11 & n_146) | (mul_68_11_n_8 & n_162));
 assign mul_68_11_n_87 = ~((n_162 | mul_68_11_n_17) & (n_152 | mul_68_11_n_11));
 assign mul_68_11_n_86 = ~((mul_68_11_n_11 & n_147) | (mul_68_11_n_16 & n_162));
 assign mul_68_11_n_85 = ~((mul_68_11_n_11 & n_148) | (mul_68_11_n_9 & n_162));
 assign mul_68_11_n_84 = ~((mul_68_11_n_11 & n_149) | (mul_68_11_n_19 & n_162));
 assign mul_68_11_n_83 = ~((mul_68_11_n_11 & n_151) | (mul_68_11_n_10 & n_162));
 assign mul_68_11_n_82 = ~((mul_68_11_n_11 & n_144) | (mul_68_11_n_15 & n_162));
 assign mul_68_11_n_81 = ~((mul_68_11_n_11 & n_150) | (mul_68_11_n_18 & n_162));
 assign mul_68_11_n_80 = ~((mul_68_11_n_11 & n_145) | (mul_68_11_n_14 & n_162));
 assign mul_68_11_n_79 = ~((mul_68_11_n_4 & n_146) | (mul_68_11_n_8 & n_154));
 assign mul_68_11_n_78 = ~((mul_68_11_n_4 & n_151) | (mul_68_11_n_10 & n_154));
 assign mul_68_11_n_77 = ~((mul_68_11_n_4 & n_152) | (mul_68_11_n_17 & n_154));
 assign mul_68_11_n_76 = ~((mul_68_11_n_4 & n_150) | (mul_68_11_n_18 & n_154));
 assign mul_68_11_n_75 = ~((n_154 | mul_68_11_n_15) & (n_144 | mul_68_11_n_4));
 assign mul_68_11_n_74 = ~((mul_68_11_n_4 & n_149) | (mul_68_11_n_19 & n_154));
 assign mul_68_11_n_73 = ~((mul_68_11_n_4 & n_145) | (mul_68_11_n_14 & n_154));
 assign mul_68_11_n_72 = ~((mul_68_11_n_4 & n_147) | (mul_68_11_n_16 & n_154));
 assign mul_68_11_n_71 = ~(n_161 ^ n_162);
 assign mul_68_11_n_70 = ((mul_68_11_n_6 & ~n_157) | (n_158 & n_157));
 assign mul_68_11_n_69 = ~(n_156 ^ n_155);
 assign mul_68_11_n_68 = ~(n_159 ^ n_160);
 assign mul_68_11_n_58 = ~mul_68_11_n_57;
 assign mul_68_11_n_39 = ~mul_68_11_n_38;
 assign mul_68_11_n_37 = ~((mul_68_11_n_12 & n_153) | (mul_68_11_n_7 & n_156));
 assign mul_68_11_n_36 = ~((mul_68_11_n_5 & n_153) | (mul_68_11_n_7 & n_160));
 assign mul_68_11_n_35 = ~((mul_68_11_n_6 & n_153) | (mul_68_11_n_7 & n_158));
 assign mul_68_11_n_34 = ~((mul_68_11_n_4 & n_153) | (mul_68_11_n_7 & n_154));
 assign mul_68_11_n_33 = ~((n_162 | mul_68_11_n_7) & (n_153 | mul_68_11_n_11));
 assign mul_68_11_n_32 = ~((n_163 | mul_68_11_n_11) & (n_162 | mul_68_11_n_13));
 assign mul_68_11_n_63 = ~((mul_68_11_n_12 & n_152) | (mul_68_11_n_17 & n_156));
 assign mul_68_11_n_62 = ~((mul_68_11_n_6 & n_151) | (mul_68_11_n_10 & n_158));
 assign mul_68_11_n_61 = ~((mul_68_11_n_5 & n_149) | (mul_68_11_n_19 & n_160));
 assign mul_68_11_n_60 = ~((mul_68_11_n_12 & n_149) | (mul_68_11_n_19 & n_156));
 assign mul_68_11_n_59 = ~((mul_68_11_n_6 & n_147) | (mul_68_11_n_16 & n_158));
 assign mul_68_11_n_57 = ~((mul_68_11_n_12 & n_144) | (mul_68_11_n_15 & n_156));
 assign mul_68_11_n_56 = ~((mul_68_11_n_12 & n_147) | (mul_68_11_n_16 & n_156));
 assign mul_68_11_n_55 = ~((mul_68_11_n_5 & n_151) | (mul_68_11_n_10 & n_160));
 assign mul_68_11_n_54 = ~((mul_68_11_n_12 & n_146) | (mul_68_11_n_8 & n_156));
 assign mul_68_11_n_53 = ~((mul_68_11_n_6 & n_146) | (mul_68_11_n_8 & n_158));
 assign mul_68_11_n_52 = ~((mul_68_11_n_6 & n_149) | (mul_68_11_n_19 & n_158));
 assign mul_68_11_n_51 = ~((mul_68_11_n_6 & n_152) | (mul_68_11_n_17 & n_158));
 assign mul_68_11_n_50 = ~((mul_68_11_n_12 & n_148) | (mul_68_11_n_9 & n_156));
 assign mul_68_11_n_49 = ~((mul_68_11_n_5 & n_145) | (mul_68_11_n_14 & n_160));
 assign mul_68_11_n_48 = ~((mul_68_11_n_5 & n_146) | (mul_68_11_n_8 & n_160));
 assign mul_68_11_n_47 = ~((mul_68_11_n_6 & n_145) | (mul_68_11_n_14 & n_158));
 assign mul_68_11_n_46 = ~((mul_68_11_n_12 & n_150) | (mul_68_11_n_18 & n_156));
 assign mul_68_11_n_45 = ~((mul_68_11_n_12 & n_151) | (mul_68_11_n_10 & n_156));
 assign mul_68_11_n_44 = ~((mul_68_11_n_6 & n_150) | (mul_68_11_n_18 & n_158));
 assign mul_68_11_n_43 = ~((mul_68_11_n_12 & n_145) | (mul_68_11_n_14 & n_156));
 assign mul_68_11_n_42 = ~((mul_68_11_n_5 & n_148) | (mul_68_11_n_9 & n_160));
 assign mul_68_11_n_41 = ~((mul_68_11_n_5 & n_152) | (mul_68_11_n_17 & n_160));
 assign mul_68_11_n_40 = ~((mul_68_11_n_6 & n_148) | (mul_68_11_n_9 & n_158));
 assign mul_68_11_n_38 = ~((mul_68_11_n_5 & n_144) | (mul_68_11_n_15 & n_160));
 assign mul_68_11_n_29 = ~(mul_68_11_n_4 | mul_68_11_n_18);
 assign mul_68_11_n_28 = ~(mul_68_11_n_4 | mul_68_11_n_17);
 assign mul_68_11_n_30 = ~(n_154 & n_147);
 assign mul_68_11_n_25 = ~(mul_68_11_n_5 & mul_68_11_n_7);
 assign mul_68_11_n_24 = ~(n_154 & n_144);
 assign mul_68_11_n_23 = ~(mul_68_11_n_4 | mul_68_11_n_10);
 assign mul_68_11_n_22 = ~(mul_68_11_n_4 | mul_68_11_n_8);
 assign mul_68_11_n_21 = ~(mul_68_11_n_4 | mul_68_11_n_7);
 assign mul_68_11_n_20 = ~(mul_68_11_n_4 | mul_68_11_n_9);
 assign mul_68_11_n_27 = ~(n_154 & n_145);
 assign mul_68_11_n_26 = ~(n_154 & n_149);
 assign mul_68_11_n_19 = ~n_149;
 assign mul_68_11_n_18 = ~n_150;
 assign mul_68_11_n_17 = ~n_152;
 assign mul_68_11_n_16 = ~n_147;
 assign mul_68_11_n_15 = ~n_144;
 assign mul_68_11_n_14 = ~n_145;
 assign mul_68_11_n_13 = ~n_163;
 assign mul_68_11_n_12 = ~n_156;
 assign mul_68_11_n_11 = ~n_162;
 assign mul_68_11_n_10 = ~n_151;
 assign mul_68_11_n_9 = ~n_148;
 assign mul_68_11_n_8 = ~n_146;
 assign mul_68_11_n_7 = ~n_153;
 assign mul_68_11_n_6 = ~n_158;
 assign mul_68_11_n_5 = ~n_160;
 assign mul_68_11_n_4 = ~n_154;
 assign mul_68_11_n_2 = ~(mul_68_11_n_12 & ~n_155);
 assign mul_68_11_n_1 = ~(mul_68_11_n_6 & ~n_157);
 assign mul_68_11_n_0 = ~(mul_68_11_n_11 & ~n_161);
 assign mul_71_11_n_5 = (mul_71_11_n_138 | (mul_71_11_n_139 & mul_71_11_n_99));
 assign {out1[28]} = ~(mul_71_11_n_541 ^ mul_71_11_n_305);
 assign {out1[27]} = ~(mul_71_11_n_542 ^ mul_71_11_n_348);
 assign {out1[23]} = ~(mul_71_11_n_537 ^ mul_71_11_n_441);
 assign mul_71_11_n_542 = ~(mul_71_11_n_358 & (mul_71_11_n_534 | mul_71_11_n_353));
 assign mul_71_11_n_541 = ~(mul_71_11_n_455 & (mul_71_11_n_538 & (mul_71_11_n_358 | mul_71_11_n_344)));
 assign {out1[26]} = ~(mul_71_11_n_534 ^ mul_71_11_n_366);
 assign {out1[25]} = ~(mul_71_11_n_533 ^ mul_71_11_n_389);
 assign mul_71_11_n_538 = ~(mul_71_11_n_329 | (mul_71_11_n_525 & (mul_71_11_n_411 & mul_71_11_n_365)));
 assign mul_71_11_n_537 = ~(mul_71_11_n_415 & (mul_71_11_n_530 | mul_71_11_n_416));
 assign {out1[22]} = ~(mul_71_11_n_530 ^ mul_71_11_n_442);
 assign {out1[21]} = ~(mul_71_11_n_529 ^ mul_71_11_n_443);
 assign mul_71_11_n_534 = ~(mul_71_11_n_439 | (mul_71_11_n_525 & mul_71_11_n_411));
 assign mul_71_11_n_533 = ~(mul_71_11_n_390 & (mul_71_11_n_526 | mul_71_11_n_388));
 assign {out1[24]} = ~(mul_71_11_n_526 ^ mul_71_11_n_412);
 assign {out1[19]} = ~(mul_71_11_n_527 ^ mul_71_11_n_430);
 assign mul_71_11_n_530 = ~(mul_71_11_n_457 | (mul_71_11_n_438 & mul_71_11_n_522));
 assign mul_71_11_n_529 = ~(mul_71_11_n_407 & ~(mul_71_11_n_522 & mul_71_11_n_406));
 assign {out1[20]} = ~(mul_71_11_n_522 ^ mul_71_11_n_444);
 assign mul_71_11_n_527 = ~(mul_71_11_n_449 & (mul_71_11_n_519 | mul_71_11_n_446));
 assign mul_71_11_n_526 = ~mul_71_11_n_525;
 assign mul_71_11_n_525 = ~(mul_71_11_n_504 & (mul_71_11_n_520 | mul_71_11_n_458));
 assign {out1[18]} = ~(mul_71_11_n_519 ^ mul_71_11_n_464);
 assign {out1[17]} = ~(mul_71_11_n_518 ^ mul_71_11_n_463);
 assign mul_71_11_n_522 = ~(mul_71_11_n_520 & ~mul_71_11_n_492);
 assign {out1[15]} = ~(mul_71_11_n_516 ^ mul_71_11_n_461);
 assign mul_71_11_n_520 = ~(mul_71_11_n_515 & mul_71_11_n_466);
 assign mul_71_11_n_519 = ~(mul_71_11_n_515 | mul_71_11_n_473);
 assign mul_71_11_n_518 = ~(mul_71_11_n_448 & (mul_71_11_n_512 | mul_71_11_n_437));
 assign {out1[16]} = ~(mul_71_11_n_512 ^ mul_71_11_n_462);
 assign mul_71_11_n_516 = ~(mul_71_11_n_447 & (mul_71_11_n_434 | mul_71_11_n_511));
 assign mul_71_11_n_515 = ~(mul_71_11_n_435 | (mul_71_11_n_437 | mul_71_11_n_512));
 assign {out1[14]} = ~(mul_71_11_n_511 ^ mul_71_11_n_453);
 assign {out1[13]} = ~(mul_71_11_n_510 ^ mul_71_11_n_429);
 assign mul_71_11_n_512 = ~(mul_71_11_n_509 | ~(mul_71_11_n_498 | mul_71_11_n_496));
 assign mul_71_11_n_511 = ~(mul_71_11_n_494 | (mul_71_11_n_506 & mul_71_11_n_485));
 assign mul_71_11_n_510 = ~(mul_71_11_n_479 & ~(mul_71_11_n_506 & mul_71_11_n_475));
 assign mul_71_11_n_509 = ~(mul_71_11_n_452 & (mul_71_11_n_501 & (mul_71_11_n_500 | mul_71_11_n_496)));
 assign {out1[12]} = ~(mul_71_11_n_506 ^ mul_71_11_n_488);
 assign {out1[11]} = ~(mul_71_11_n_505 ^ mul_71_11_n_487);
 assign mul_71_11_n_506 = ~(mul_71_11_n_500 & mul_71_11_n_498);
 assign mul_71_11_n_505 = ~(mul_71_11_n_477 & (mul_71_11_n_499 | mul_71_11_n_481));
 assign mul_71_11_n_504 = ~(mul_71_11_n_433 | (mul_71_11_n_502 | (mul_71_11_n_457 & mul_71_11_n_440)));
 assign {out1[10]} = ~(mul_71_11_n_489 ^ mul_71_11_n_499);
 assign mul_71_11_n_502 = ~(mul_71_11_n_410 & ~(mul_71_11_n_492 & mul_71_11_n_459));
 assign mul_71_11_n_501 = ~(mul_71_11_n_465 | (mul_71_11_n_494 & mul_71_11_n_460));
 assign mul_71_11_n_500 = ~(mul_71_11_n_490 | (mul_71_11_n_478 | (mul_71_11_n_493 & mul_71_11_n_484)));
 assign mul_71_11_n_499 = ~(mul_71_11_n_495 | mul_71_11_n_493);
 assign mul_71_11_n_498 = ~(mul_71_11_n_495 & mul_71_11_n_484);
 assign {out1[9]} = ~(mul_71_11_n_483 ^ mul_71_11_n_486);
 assign mul_71_11_n_496 = ~(mul_71_11_n_460 & mul_71_11_n_485);
 assign mul_71_11_n_495 = ~(mul_71_11_n_480 | (mul_71_11_n_445 | mul_71_11_n_456));
 assign mul_71_11_n_494 = ~(mul_71_11_n_418 & (mul_71_11_n_479 | mul_71_11_n_414));
 assign mul_71_11_n_493 = ~(mul_71_11_n_476 & (mul_71_11_n_480 | mul_71_11_n_450));
 assign mul_71_11_n_492 = ~(mul_71_11_n_409 & (mul_71_11_n_491 & (mul_71_11_n_449 | mul_71_11_n_413)));
 assign mul_71_11_n_491 = ~(mul_71_11_n_473 & mul_71_11_n_466);
 assign mul_71_11_n_490 = ~(mul_71_11_n_477 | mul_71_11_n_474);
 assign mul_71_11_n_489 = ~(mul_71_11_n_481 | ~mul_71_11_n_477);
 assign mul_71_11_n_488 = ~(mul_71_11_n_475 & mul_71_11_n_479);
 assign mul_71_11_n_487 = (mul_71_11_n_474 | mul_71_11_n_478);
 assign mul_71_11_n_486 = ~(mul_71_11_n_476 & ~mul_71_11_n_480);
 assign mul_71_11_n_485 = ~(mul_71_11_n_414 | ~mul_71_11_n_475);
 assign mul_71_11_n_484 = ~(mul_71_11_n_481 | mul_71_11_n_474);
 assign mul_71_11_n_483 = ~(mul_71_11_n_450 & (mul_71_11_n_456 | mul_71_11_n_445));
 assign {out1[8]} = ~(mul_71_11_n_456 ^ mul_71_11_n_454);
 assign mul_71_11_n_481 = ~(mul_71_11_n_470 | mul_71_11_n_467);
 assign mul_71_11_n_480 = ~(mul_71_11_n_468 | mul_71_11_n_419);
 assign mul_71_11_n_479 = ~(mul_71_11_n_401 & mul_71_11_n_471);
 assign mul_71_11_n_478 = (mul_71_11_n_472 & mul_71_11_n_469);
 assign mul_71_11_n_477 = ~(mul_71_11_n_470 & mul_71_11_n_467);
 assign mul_71_11_n_476 = ~(mul_71_11_n_468 & mul_71_11_n_419);
 assign mul_71_11_n_475 = (mul_71_11_n_401 | mul_71_11_n_471);
 assign mul_71_11_n_474 = ~(mul_71_11_n_472 | mul_71_11_n_469);
 assign mul_71_11_n_473 = ~(mul_71_11_n_451 & (mul_71_11_n_435 | mul_71_11_n_448));
 assign mul_71_11_n_471 = ((mul_71_11_n_369 & mul_71_11_n_324) | ((mul_71_11_n_324 & mul_71_11_n_275)
    | (mul_71_11_n_275 & mul_71_11_n_369)));
 assign mul_71_11_n_472 = (mul_71_11_n_324 ^ (mul_71_11_n_275 ^ mul_71_11_n_369));
 assign mul_71_11_n_469 = ((mul_71_11_n_367 & mul_71_11_n_370) | ((mul_71_11_n_370 & mul_71_11_n_285)
    | (mul_71_11_n_285 & mul_71_11_n_367)));
 assign mul_71_11_n_470 = (mul_71_11_n_370 ^ (mul_71_11_n_285 ^ mul_71_11_n_367));
 assign mul_71_11_n_467 = ((mul_71_11_n_368 & mul_71_11_n_229) | ((mul_71_11_n_229 & mul_71_11_n_356)
    | (mul_71_11_n_356 & mul_71_11_n_368)));
 assign mul_71_11_n_468 = (mul_71_11_n_229 ^ (mul_71_11_n_356 ^ mul_71_11_n_368));
 assign mul_71_11_n_465 = ~(mul_71_11_n_447 | mul_71_11_n_436);
 assign mul_71_11_n_466 = ~(mul_71_11_n_446 | mul_71_11_n_413);
 assign mul_71_11_n_464 = ~(mul_71_11_n_446 | ~mul_71_11_n_449);
 assign mul_71_11_n_463 = ~(mul_71_11_n_451 & ~mul_71_11_n_435);
 assign mul_71_11_n_462 = ~(mul_71_11_n_437 | ~mul_71_11_n_448);
 assign mul_71_11_n_461 = ~(mul_71_11_n_452 & ~mul_71_11_n_436);
 assign mul_71_11_n_459 = ~mul_71_11_n_458;
 assign mul_71_11_n_455 = ~(mul_71_11_n_439 & mul_71_11_n_365);
 assign mul_71_11_n_454 = ~(mul_71_11_n_445 | ~mul_71_11_n_450);
 assign mul_71_11_n_460 = ~(mul_71_11_n_434 | mul_71_11_n_436);
 assign mul_71_11_n_458 = ~(mul_71_11_n_438 & mul_71_11_n_440);
 assign mul_71_11_n_457 = ~(mul_71_11_n_417 & (mul_71_11_n_408 | mul_71_11_n_407));
 assign mul_71_11_n_453 = ~(mul_71_11_n_434 | ~mul_71_11_n_447);
 assign mul_71_11_n_456 = ~(mul_71_11_n_432 | ((mul_71_11_n_382 & mul_71_11_n_362) | (mul_71_11_n_391
    & mul_71_11_n_354)));
 assign mul_71_11_n_452 = ~(mul_71_11_n_426 & mul_71_11_n_421);
 assign mul_71_11_n_444 = ~(mul_71_11_n_406 & mul_71_11_n_407);
 assign mul_71_11_n_443 = ~(mul_71_11_n_417 & ~mul_71_11_n_408);
 assign mul_71_11_n_451 = ~(mul_71_11_n_428 & mul_71_11_n_423);
 assign mul_71_11_n_442 = ~(mul_71_11_n_416 | ~mul_71_11_n_415);
 assign mul_71_11_n_441 = ~(mul_71_11_n_410 & ~mul_71_11_n_405);
 assign mul_71_11_n_450 = ~(mul_71_11_n_420 & mul_71_11_n_372);
 assign mul_71_11_n_449 = ~(mul_71_11_n_395 & mul_71_11_n_427);
 assign mul_71_11_n_448 = ~(mul_71_11_n_424 & mul_71_11_n_425);
 assign mul_71_11_n_447 = ~(mul_71_11_n_422 & mul_71_11_n_396);
 assign mul_71_11_n_446 = ~(mul_71_11_n_395 | mul_71_11_n_427);
 assign mul_71_11_n_445 = ~(mul_71_11_n_420 | mul_71_11_n_372);
 assign mul_71_11_n_433 = ~(mul_71_11_n_415 | mul_71_11_n_405);
 assign mul_71_11_n_432 = ~(mul_71_11_n_383 & ~(mul_71_11_n_391 & mul_71_11_n_359));
 assign {out1[7]} = ~(mul_71_11_n_387 ^ mul_71_11_n_386);
 assign mul_71_11_n_440 = ~(mul_71_11_n_416 | mul_71_11_n_405);
 assign mul_71_11_n_430 = ~(mul_71_11_n_409 & ~mul_71_11_n_413);
 assign mul_71_11_n_429 = ~(mul_71_11_n_418 & ~mul_71_11_n_414);
 assign mul_71_11_n_439 = ~(mul_71_11_n_379 & (mul_71_11_n_390 | mul_71_11_n_380));
 assign mul_71_11_n_438 = ~(mul_71_11_n_408 | ~mul_71_11_n_406);
 assign mul_71_11_n_437 = ~(mul_71_11_n_424 | mul_71_11_n_425);
 assign mul_71_11_n_436 = ~(mul_71_11_n_426 | mul_71_11_n_421);
 assign mul_71_11_n_435 = ~(mul_71_11_n_428 | mul_71_11_n_423);
 assign mul_71_11_n_434 = ~(mul_71_11_n_422 | mul_71_11_n_396);
 assign mul_71_11_n_427 = ((mul_71_11_n_314 & mul_71_11_n_268) | ((mul_71_11_n_268 & mul_71_11_n_332)
    | (mul_71_11_n_332 & mul_71_11_n_314)));
 assign mul_71_11_n_428 = (mul_71_11_n_268 ^ (mul_71_11_n_332 ^ mul_71_11_n_314));
 assign mul_71_11_n_425 = ((mul_71_11_n_343 & mul_71_11_n_340) | ((mul_71_11_n_340 & mul_71_11_n_296)
    | (mul_71_11_n_296 & mul_71_11_n_343)));
 assign mul_71_11_n_426 = (mul_71_11_n_340 ^ (mul_71_11_n_296 ^ mul_71_11_n_343));
 assign mul_71_11_n_423 = ((mul_71_11_n_333 & mul_71_11_n_342) | ((mul_71_11_n_342 & mul_71_11_n_269)
    | (mul_71_11_n_269 & mul_71_11_n_333)));
 assign mul_71_11_n_424 = (mul_71_11_n_342 ^ (mul_71_11_n_269 ^ mul_71_11_n_333));
 assign mul_71_11_n_421 = ((mul_71_11_n_336 & mul_71_11_n_341) | ((mul_71_11_n_341 & mul_71_11_n_292)
    | (mul_71_11_n_292 & mul_71_11_n_336)));
 assign mul_71_11_n_422 = (mul_71_11_n_341 ^ (mul_71_11_n_292 ^ mul_71_11_n_336));
 assign mul_71_11_n_419 = ((mul_71_11_n_357 & mul_71_11_n_245) | ((mul_71_11_n_245 & mul_71_11_n_334)
    | (mul_71_11_n_334 & mul_71_11_n_357)));
 assign mul_71_11_n_420 = (mul_71_11_n_245 ^ (mul_71_11_n_334 ^ mul_71_11_n_357));
 assign mul_71_11_n_418 = ~(mul_71_11_n_397 & mul_71_11_n_400);
 assign mul_71_11_n_412 = ~(mul_71_11_n_388 | ~mul_71_11_n_390);
 assign mul_71_11_n_417 = ~(mul_71_11_n_377 & mul_71_11_n_402);
 assign mul_71_11_n_416 = ~(mul_71_11_n_399 | mul_71_11_n_376);
 assign mul_71_11_n_415 = ~(mul_71_11_n_399 & mul_71_11_n_376);
 assign mul_71_11_n_414 = ~(mul_71_11_n_397 | mul_71_11_n_400);
 assign mul_71_11_n_413 = ~(mul_71_11_n_393 | mul_71_11_n_394);
 assign {out1[6]} = ~(mul_71_11_n_364 ^ mul_71_11_n_381);
 assign mul_71_11_n_411 = ~(mul_71_11_n_388 | mul_71_11_n_380);
 assign mul_71_11_n_410 = ~(mul_71_11_n_385 & mul_71_11_n_398);
 assign mul_71_11_n_409 = ~(mul_71_11_n_393 & mul_71_11_n_394);
 assign mul_71_11_n_408 = ~(mul_71_11_n_377 | mul_71_11_n_402);
 assign mul_71_11_n_407 = ~(mul_71_11_n_403 & mul_71_11_n_392);
 assign mul_71_11_n_406 = (mul_71_11_n_403 | mul_71_11_n_392);
 assign mul_71_11_n_405 = ~(mul_71_11_n_385 | mul_71_11_n_398);
 assign mul_71_11_n_402 = ((mul_71_11_n_326 & mul_71_11_n_280) | ((mul_71_11_n_280 & mul_71_11_n_321)
    | (mul_71_11_n_321 & mul_71_11_n_326)));
 assign mul_71_11_n_403 = (mul_71_11_n_280 ^ (mul_71_11_n_321 ^ mul_71_11_n_326));
 assign mul_71_11_n_400 = ((mul_71_11_n_320 & mul_71_11_n_323) | ((mul_71_11_n_323 & mul_71_11_n_273)
    | (mul_71_11_n_273 & mul_71_11_n_320)));
 assign mul_71_11_n_401 = (mul_71_11_n_323 ^ (mul_71_11_n_273 ^ mul_71_11_n_320));
 assign mul_71_11_n_398 = ((mul_71_11_n_309 & mul_71_11_n_318) | ((mul_71_11_n_318 & mul_71_11_n_263)
    | (mul_71_11_n_263 & mul_71_11_n_309)));
 assign mul_71_11_n_399 = (mul_71_11_n_318 ^ (mul_71_11_n_263 ^ mul_71_11_n_309));
 assign mul_71_11_n_396 = ((mul_71_11_n_337 & mul_71_11_n_272) | ((mul_71_11_n_272 & mul_71_11_n_319)
    | (mul_71_11_n_319 & mul_71_11_n_337)));
 assign mul_71_11_n_397 = (mul_71_11_n_272 ^ (mul_71_11_n_319 ^ mul_71_11_n_337));
 assign mul_71_11_n_394 = ((mul_71_11_n_313 & mul_71_11_n_316) | ((mul_71_11_n_316 & mul_71_11_n_277)
    | (mul_71_11_n_277 & mul_71_11_n_313)));
 assign mul_71_11_n_395 = (mul_71_11_n_316 ^ (mul_71_11_n_277 ^ mul_71_11_n_313));
 assign mul_71_11_n_392 = ((mul_71_11_n_322 & mul_71_11_n_315) | ((mul_71_11_n_315 & mul_71_11_n_281)
    | (mul_71_11_n_281 & mul_71_11_n_322)));
 assign mul_71_11_n_393 = (mul_71_11_n_315 ^ (mul_71_11_n_281 ^ mul_71_11_n_322));
 assign mul_71_11_n_391 = ~(mul_71_11_n_371 | ~mul_71_11_n_382);
 assign mul_71_11_n_389 = ~(mul_71_11_n_379 & ~mul_71_11_n_380);
 assign mul_71_11_n_390 = ~(mul_71_11_n_375 & mul_71_11_n_384);
 assign mul_71_11_n_387 = ~(mul_71_11_n_382 & mul_71_11_n_383);
 assign mul_71_11_n_386 = ~(mul_71_11_n_363 & (mul_71_11_n_364 | mul_71_11_n_371));
 assign mul_71_11_n_388 = ~(mul_71_11_n_375 | mul_71_11_n_384);
 assign mul_71_11_n_384 = ((mul_71_11_n_317 & mul_71_11_n_308) | ((mul_71_11_n_308 & mul_71_11_n_278)
    | (mul_71_11_n_278 & mul_71_11_n_317)));
 assign mul_71_11_n_385 = (mul_71_11_n_308 ^ (mul_71_11_n_278 ^ mul_71_11_n_317));
 assign mul_71_11_n_383 = ~(mul_71_11_n_373 & mul_71_11_n_360);
 assign mul_71_11_n_382 = (mul_71_11_n_373 | mul_71_11_n_360);
 assign mul_71_11_n_381 = ~(mul_71_11_n_371 | mul_71_11_n_362);
 assign mul_71_11_n_380 = ~(mul_71_11_n_351 | mul_71_11_n_374);
 assign mul_71_11_n_379 = ~(mul_71_11_n_351 & mul_71_11_n_374);
 assign {out1[5]} = ~(mul_71_11_n_347 ^ mul_71_11_n_355);
 assign mul_71_11_n_376 = ((mul_71_11_n_310 & mul_71_11_n_265) | ((mul_71_11_n_265 & mul_71_11_n_325)
    | (mul_71_11_n_325 & mul_71_11_n_310)));
 assign mul_71_11_n_377 = (mul_71_11_n_265 ^ (mul_71_11_n_325 ^ mul_71_11_n_310));
 assign mul_71_11_n_374 = ((mul_71_11_n_307 & mul_71_11_n_261) | ((mul_71_11_n_261 & mul_71_11_n_302)
    | (mul_71_11_n_302 & mul_71_11_n_307)));
 assign mul_71_11_n_375 = (mul_71_11_n_261 ^ (mul_71_11_n_302 ^ mul_71_11_n_307));
 assign mul_71_11_n_369 = ((mul_71_11_n_338 & mul_71_11_n_243) | ((mul_71_11_n_243 & mul_71_11_n_150)
    | (mul_71_11_n_150 & mul_71_11_n_338)));
 assign mul_71_11_n_370 = (mul_71_11_n_243 ^ (mul_71_11_n_150 ^ mul_71_11_n_338));
 assign mul_71_11_n_367 = ((mul_71_11_n_339 & mul_71_11_n_165) | ((mul_71_11_n_165 & mul_71_11_n_208)
    | (mul_71_11_n_208 & mul_71_11_n_339)));
 assign mul_71_11_n_368 = (mul_71_11_n_165 ^ (mul_71_11_n_208 ^ mul_71_11_n_339));
 assign mul_71_11_n_372 = ((mul_71_11_n_335 & mul_71_11_n_228) | ((mul_71_11_n_228 & mul_71_11_n_162)
    | (mul_71_11_n_162 & mul_71_11_n_335)));
 assign mul_71_11_n_373 = (mul_71_11_n_228 ^ (mul_71_11_n_162 ^ mul_71_11_n_335));
 assign mul_71_11_n_366 = ~(mul_71_11_n_353 | ~mul_71_11_n_358);
 assign mul_71_11_n_371 = ~(mul_71_11_n_361 | mul_71_11_n_311);
 assign mul_71_11_n_363 = ~mul_71_11_n_362;
 assign mul_71_11_n_365 = ~(mul_71_11_n_353 | mul_71_11_n_344);
 assign mul_71_11_n_364 = ~(mul_71_11_n_354 | mul_71_11_n_359);
 assign mul_71_11_n_362 = (mul_71_11_n_361 & mul_71_11_n_311);
 assign mul_71_11_n_356 = ((mul_71_11_n_300 & mul_71_11_n_159) | ((mul_71_11_n_159 & mul_71_11_n_207)
    | (mul_71_11_n_207 & mul_71_11_n_300)));
 assign mul_71_11_n_357 = (mul_71_11_n_159 ^ (mul_71_11_n_207 ^ mul_71_11_n_300));
 assign mul_71_11_n_360 = ((mul_71_11_n_298 & mul_71_11_n_230) | ((mul_71_11_n_230 & mul_71_11_n_160)
    | (mul_71_11_n_160 & mul_71_11_n_298)));
 assign mul_71_11_n_361 = (mul_71_11_n_230 ^ (mul_71_11_n_160 ^ mul_71_11_n_298));
 assign mul_71_11_n_359 = ~(mul_71_11_n_345 | mul_71_11_n_349);
 assign mul_71_11_n_355 = ~(mul_71_11_n_349 & mul_71_11_n_289);
 assign mul_71_11_n_358 = ~(mul_71_11_n_350 & mul_71_11_n_328);
 assign {out1[4]} = ~(mul_71_11_n_306 ^ mul_71_11_n_346);
 assign mul_71_11_n_354 = ~(mul_71_11_n_330 & (mul_71_11_n_345 | mul_71_11_n_289));
 assign mul_71_11_n_353 = ~(mul_71_11_n_350 | mul_71_11_n_328);
 assign mul_71_11_n_350 = ((mul_71_11_n_283 & mul_71_11_n_301) | ((mul_71_11_n_301 & mul_71_11_n_189)
    | (mul_71_11_n_189 & mul_71_11_n_283)));
 assign mul_71_11_n_351 = (mul_71_11_n_301 ^ (mul_71_11_n_189 ^ mul_71_11_n_283));
 assign mul_71_11_n_349 = ~(mul_71_11_n_346 & mul_71_11_n_290);
 assign mul_71_11_n_348 = (mul_71_11_n_344 | mul_71_11_n_329);
 assign mul_71_11_n_347 = ~(mul_71_11_n_330 & ~mul_71_11_n_345);
 assign mul_71_11_n_342 = ((mul_71_11_n_291 & mul_71_11_n_246) | ((mul_71_11_n_246 & mul_71_11_n_157)
    | (mul_71_11_n_157 & mul_71_11_n_291)));
 assign mul_71_11_n_343 = (mul_71_11_n_246 ^ (mul_71_11_n_157 ^ mul_71_11_n_291));
 assign mul_71_11_n_340 = ((mul_71_11_n_303 & mul_71_11_n_231) | ((mul_71_11_n_231 & mul_71_11_n_151)
    | (mul_71_11_n_151 & mul_71_11_n_303)));
 assign mul_71_11_n_341 = (mul_71_11_n_231 ^ (mul_71_11_n_151 ^ mul_71_11_n_303));
 assign mul_71_11_n_338 = ((mul_71_11_n_299 & mul_71_11_n_203) | ((mul_71_11_n_203 & mul_71_11_n_149)
    | (mul_71_11_n_149 & mul_71_11_n_299)));
 assign mul_71_11_n_339 = (mul_71_11_n_203 ^ (mul_71_11_n_149 ^ mul_71_11_n_299));
 assign mul_71_11_n_336 = ((mul_71_11_n_304 & mul_71_11_n_234) | ((mul_71_11_n_234 & mul_71_11_n_166)
    | (mul_71_11_n_166 & mul_71_11_n_304)));
 assign mul_71_11_n_337 = (mul_71_11_n_234 ^ (mul_71_11_n_166 ^ mul_71_11_n_304));
 assign mul_71_11_n_334 = ((mul_71_11_n_297 & mul_71_11_n_202) | ((mul_71_11_n_202 & mul_71_11_n_258)
    | (mul_71_11_n_258 & mul_71_11_n_297)));
 assign mul_71_11_n_335 = (mul_71_11_n_202 ^ (mul_71_11_n_258 ^ mul_71_11_n_297));
 assign mul_71_11_n_332 = ((mul_71_11_n_295 & mul_71_11_n_244) | ((mul_71_11_n_244 & mul_71_11_n_161)
    | (mul_71_11_n_161 & mul_71_11_n_295)));
 assign mul_71_11_n_333 = (mul_71_11_n_244 ^ (mul_71_11_n_161 ^ mul_71_11_n_295));
 assign mul_71_11_n_346 = ((mul_71_11_n_293 & mul_71_11_n_249) | ((mul_71_11_n_249 & mul_71_11_n_256)
    | (mul_71_11_n_256 & mul_71_11_n_293)));
 assign {out1[3]} = (mul_71_11_n_249 ^ (mul_71_11_n_256 ^ mul_71_11_n_293));
 assign mul_71_11_n_345 = ~(mul_71_11_n_312 | mul_71_11_n_287);
 assign mul_71_11_n_344 = ~(mul_71_11_n_327 | mul_71_11_n_286);
 assign mul_71_11_n_330 = ~(mul_71_11_n_312 & mul_71_11_n_287);
 assign mul_71_11_n_329 = (mul_71_11_n_327 & mul_71_11_n_286);
 assign mul_71_11_n_327 = ((mul_71_11_n_282 & mul_71_11_n_186) | ((mul_71_11_n_186 & mul_71_11_n_242)
    | (mul_71_11_n_242 & mul_71_11_n_282)));
 assign mul_71_11_n_328 = (mul_71_11_n_186 ^ (mul_71_11_n_242 ^ mul_71_11_n_282));
 assign mul_71_11_n_325 = ((mul_71_11_n_266 & mul_71_11_n_232) | ((mul_71_11_n_232 & mul_71_11_n_156)
    | (mul_71_11_n_156 & mul_71_11_n_266)));
 assign mul_71_11_n_326 = (mul_71_11_n_232 ^ (mul_71_11_n_156 ^ mul_71_11_n_266));
 assign mul_71_11_n_323 = ((mul_71_11_n_284 & mul_71_11_n_238) | ((mul_71_11_n_238 & mul_71_11_n_154)
    | (mul_71_11_n_154 & mul_71_11_n_284)));
 assign mul_71_11_n_324 = (mul_71_11_n_238 ^ (mul_71_11_n_154 ^ mul_71_11_n_284));
 assign mul_71_11_n_321 = ((mul_71_11_n_276 & mul_71_11_n_240) | ((mul_71_11_n_240 & mul_71_11_n_153)
    | (mul_71_11_n_153 & mul_71_11_n_276)));
 assign mul_71_11_n_322 = (mul_71_11_n_240 ^ (mul_71_11_n_153 ^ mul_71_11_n_276));
 assign mul_71_11_n_319 = ((mul_71_11_n_274 & mul_71_11_n_235) | ((mul_71_11_n_235 & mul_71_11_n_152)
    | (mul_71_11_n_152 & mul_71_11_n_274)));
 assign mul_71_11_n_320 = (mul_71_11_n_235 ^ (mul_71_11_n_152 ^ mul_71_11_n_274));
 assign mul_71_11_n_317 = ((mul_71_11_n_279 & mul_71_11_n_3) | ((mul_71_11_n_3 & mul_71_11_n_193) | (mul_71_11_n_193
    & mul_71_11_n_279)));
 assign mul_71_11_n_318 = (mul_71_11_n_3 ^ (mul_71_11_n_193 ^ mul_71_11_n_279));
 assign mul_71_11_n_315 = ((mul_71_11_n_270 & mul_71_11_n_233) | ((mul_71_11_n_233 & mul_71_11_n_167)
    | (mul_71_11_n_167 & mul_71_11_n_270)));
 assign mul_71_11_n_316 = (mul_71_11_n_233 ^ (mul_71_11_n_167 ^ mul_71_11_n_270));
 assign mul_71_11_n_313 = ((mul_71_11_n_271 & mul_71_11_n_236) | ((mul_71_11_n_236 & mul_71_11_n_164)
    | (mul_71_11_n_164 & mul_71_11_n_271)));
 assign mul_71_11_n_314 = (mul_71_11_n_236 ^ (mul_71_11_n_164 ^ mul_71_11_n_271));
 assign mul_71_11_n_311 = ((mul_71_11_n_260 & mul_71_11_n_239) | ((mul_71_11_n_239 & mul_71_11_n_155)
    | (mul_71_11_n_155 & mul_71_11_n_260)));
 assign mul_71_11_n_312 = (mul_71_11_n_239 ^ (mul_71_11_n_155 ^ mul_71_11_n_260));
 assign mul_71_11_n_309 = ((mul_71_11_n_264 & mul_71_11_n_163) | ((mul_71_11_n_163 & mul_71_11_n_206)
    | (mul_71_11_n_206 & mul_71_11_n_264)));
 assign mul_71_11_n_310 = (mul_71_11_n_163 ^ (mul_71_11_n_206 ^ mul_71_11_n_264));
 assign mul_71_11_n_307 = ((mul_71_11_n_262 & mul_71_11_n_200) | ((mul_71_11_n_200 & mul_71_11_n_205)
    | (mul_71_11_n_205 & mul_71_11_n_262)));
 assign mul_71_11_n_308 = (mul_71_11_n_200 ^ (mul_71_11_n_205 ^ mul_71_11_n_262));
 assign mul_71_11_n_306 = ~(mul_71_11_n_290 & mul_71_11_n_289);
 assign mul_71_11_n_305 = ~(mul_71_11_n_267 ^ mul_71_11_n_148);
 assign mul_71_11_n_303 = ((mul_71_11_n_212 & mul_71_11_n_177) | ((mul_71_11_n_177 & mul_71_11_n_222)
    | (mul_71_11_n_222 & mul_71_11_n_212)));
 assign mul_71_11_n_304 = (mul_71_11_n_177 ^ (mul_71_11_n_222 ^ mul_71_11_n_212));
 assign mul_71_11_n_301 = ((mul_71_11_n_5 & mul_71_11_n_188) | ((mul_71_11_n_188 & mul_71_11_n_190) |
    (mul_71_11_n_190 & mul_71_11_n_5)));
 assign mul_71_11_n_302 = (mul_71_11_n_188 ^ (mul_71_11_n_190 ^ mul_71_11_n_5));
 assign mul_71_11_n_299 = ((mul_71_11_n_257 & mul_71_11_n_197) | ((mul_71_11_n_197 & mul_71_11_n_133)
    | (mul_71_11_n_133 & mul_71_11_n_257)));
 assign mul_71_11_n_300 = (mul_71_11_n_197 ^ (mul_71_11_n_133 ^ mul_71_11_n_257));
 assign mul_71_11_n_297 = ((mul_71_11_n_259 & mul_71_11_n_204) | ((mul_71_11_n_204 & mul_71_11_n_147)
    | (mul_71_11_n_147 & mul_71_11_n_259)));
 assign mul_71_11_n_298 = (mul_71_11_n_204 ^ (mul_71_11_n_147 ^ mul_71_11_n_259));
 assign mul_71_11_n_295 = ((mul_71_11_n_211 & mul_71_11_n_169) | ((mul_71_11_n_169 & mul_71_11_n_225)
    | (mul_71_11_n_225 & mul_71_11_n_211)));
 assign mul_71_11_n_296 = (mul_71_11_n_169 ^ (mul_71_11_n_225 ^ mul_71_11_n_211));
 assign mul_71_11_n_293 = ((mul_71_11_n_253 & mul_71_11_n_250) | ((mul_71_11_n_250 & mul_71_11_n_132)
    | (mul_71_11_n_132 & mul_71_11_n_253)));
 assign {out1[2]} = (mul_71_11_n_250 ^ (mul_71_11_n_132 ^ mul_71_11_n_253));
 assign mul_71_11_n_291 = ((mul_71_11_n_210 & mul_71_11_n_179) | ((mul_71_11_n_179 & mul_71_11_n_223)
    | (mul_71_11_n_223 & mul_71_11_n_210)));
 assign mul_71_11_n_292 = (mul_71_11_n_179 ^ (mul_71_11_n_223 ^ mul_71_11_n_210));
 assign mul_71_11_n_290 = ~(mul_71_11_n_251 & ~mul_71_11_n_288);
 assign mul_71_11_n_289 = ~(mul_71_11_n_288 & ~mul_71_11_n_251);
 assign mul_71_11_n_287 = ((mul_71_11_n_255 & mul_71_11_n_158) | ((mul_71_11_n_158 & mul_71_11_n_146)
    | (mul_71_11_n_146 & mul_71_11_n_255)));
 assign mul_71_11_n_288 = (mul_71_11_n_158 ^ (mul_71_11_n_146 ^ mul_71_11_n_255));
 assign mul_71_11_n_284 = ((mul_71_11_n_220 & mul_71_11_n_196) | ((mul_71_11_n_196 & mul_71_11_n_178)
    | (mul_71_11_n_178 & mul_71_11_n_220)));
 assign mul_71_11_n_285 = (mul_71_11_n_196 ^ (mul_71_11_n_178 ^ mul_71_11_n_220));
 assign mul_71_11_n_282 = ((mul_71_11_n_180 & mul_71_11_n_226) | ((mul_71_11_n_226 & mul_71_11_n_241)
    | (mul_71_11_n_241 & mul_71_11_n_180)));
 assign mul_71_11_n_283 = (mul_71_11_n_226 ^ (mul_71_11_n_241 ^ mul_71_11_n_180));
 assign mul_71_11_n_280 = ((mul_71_11_n_214 & mul_71_11_n_199) | ((mul_71_11_n_199 & mul_71_11_n_176)
    | (mul_71_11_n_176 & mul_71_11_n_214)));
 assign mul_71_11_n_281 = (mul_71_11_n_199 ^ (mul_71_11_n_176 ^ mul_71_11_n_214));
 assign mul_71_11_n_276 = ((mul_71_11_n_218 & mul_71_11_n_194) | ((mul_71_11_n_194 & mul_71_11_n_173)
    | (mul_71_11_n_173 & mul_71_11_n_218)));
 assign mul_71_11_n_277 = (mul_71_11_n_194 ^ (mul_71_11_n_173 ^ mul_71_11_n_218));
 assign mul_71_11_n_274 = ((mul_71_11_n_217 & mul_71_11_n_192) | ((mul_71_11_n_192 & mul_71_11_n_171)
    | (mul_71_11_n_171 & mul_71_11_n_217)));
 assign mul_71_11_n_275 = (mul_71_11_n_192 ^ (mul_71_11_n_171 ^ mul_71_11_n_217));
 assign mul_71_11_n_272 = ((mul_71_11_n_219 & mul_71_11_n_195) | ((mul_71_11_n_195 & mul_71_11_n_172)
    | (mul_71_11_n_172 & mul_71_11_n_219)));
 assign mul_71_11_n_273 = (mul_71_11_n_195 ^ (mul_71_11_n_172 ^ mul_71_11_n_219));
 assign mul_71_11_n_270 = ((mul_71_11_n_216 & mul_71_11_n_191) | ((mul_71_11_n_191 & mul_71_11_n_170)
    | (mul_71_11_n_170 & mul_71_11_n_216)));
 assign mul_71_11_n_271 = (mul_71_11_n_191 ^ (mul_71_11_n_170 ^ mul_71_11_n_216));
 assign mul_71_11_n_268 = ((mul_71_11_n_182 & mul_71_11_n_198) | ((mul_71_11_n_198 & mul_71_11_n_227)
    | (mul_71_11_n_227 & mul_71_11_n_182)));
 assign mul_71_11_n_269 = (mul_71_11_n_198 ^ (mul_71_11_n_227 ^ mul_71_11_n_182));
 assign mul_71_11_n_267 = ((mul_71_11_n_183 & mul_71_11_n_187) | ((mul_71_11_n_187 & mul_71_11_n_237)
    | (mul_71_11_n_237 & mul_71_11_n_183)));
 assign mul_71_11_n_286 = (mul_71_11_n_187 ^ (mul_71_11_n_237 ^ mul_71_11_n_183));
 assign mul_71_11_n_265 = ((mul_71_11_n_181 & mul_71_11_n_201) | ((mul_71_11_n_201 & mul_71_11_n_224)
    | (mul_71_11_n_224 & mul_71_11_n_181)));
 assign mul_71_11_n_266 = (mul_71_11_n_201 ^ (mul_71_11_n_224 ^ mul_71_11_n_181));
 assign mul_71_11_n_261 = ((mul_71_11_n_185 & mul_71_11_n_175) | ((mul_71_11_n_175 & mul_71_11_n_19)
    | (mul_71_11_n_19 & mul_71_11_n_185)));
 assign mul_71_11_n_262 = (mul_71_11_n_175 ^ (mul_71_11_n_19 ^ mul_71_11_n_185));
 assign mul_71_11_n_259 = (mul_71_11_n_213 & mul_71_11_n_248);
 assign mul_71_11_n_260 = (mul_71_11_n_213 ^ mul_71_11_n_248);
 assign mul_71_11_n_257 = (mul_71_11_n_221 & mul_71_11_n_247);
 assign mul_71_11_n_258 = (mul_71_11_n_221 ^ mul_71_11_n_247);
 assign mul_71_11_n_255 = (mul_71_11_n_168 & mul_71_11_n_137);
 assign mul_71_11_n_256 = (mul_71_11_n_168 ^ mul_71_11_n_137);
 assign {out1[1]} = ~(mul_71_11_n_253 | (mul_71_11_n_252 & mul_71_11_n_128));
 assign mul_71_11_n_253 = ~(mul_71_11_n_252 | mul_71_11_n_128);
 assign mul_71_11_n_250 = ~((mul_71_11_n_144 | mul_71_11_n_122) & (mul_71_11_n_109 | mul_71_11_n_21));
 assign mul_71_11_n_249 = ~((mul_71_11_n_144 | mul_71_11_n_109) & (mul_71_11_n_112 | mul_71_11_n_21));
 assign mul_71_11_n_246 = ~((mul_71_11_n_144 | mul_71_11_n_115) & (mul_71_11_n_117 | mul_71_11_n_21));
 assign mul_71_11_n_245 = ~((mul_71_11_n_144 | mul_71_11_n_119) & (mul_71_11_n_110 | mul_71_11_n_21));
 assign mul_71_11_n_244 = ~((mul_71_11_n_144 | mul_71_11_n_117) & (mul_71_11_n_108 | mul_71_11_n_21));
 assign mul_71_11_n_243 = ~((mul_71_11_n_144 | mul_71_11_n_105) & (mul_71_11_n_111 | mul_71_11_n_21));
 assign mul_71_11_n_242 = ~(mul_71_11_n_142 & ~(mul_71_11_n_143 & mul_71_11_n_44));
 assign mul_71_11_n_240 = ~((mul_71_11_n_144 | mul_71_11_n_123) & (mul_71_11_n_116 | mul_71_11_n_21));
 assign mul_71_11_n_239 = ~((mul_71_11_n_144 | mul_71_11_n_102) & (mul_71_11_n_120 | mul_71_11_n_21));
 assign mul_71_11_n_238 = ~((mul_71_11_n_144 | mul_71_11_n_111) & (mul_71_11_n_104 | mul_71_11_n_21));
 assign mul_71_11_n_236 = ~((mul_71_11_n_144 | mul_71_11_n_108) & (mul_71_11_n_106 | mul_71_11_n_21));
 assign mul_71_11_n_235 = ~((mul_71_11_n_144 | mul_71_11_n_104) & (mul_71_11_n_107 | mul_71_11_n_21));
 assign mul_71_11_n_234 = ~((mul_71_11_n_144 | mul_71_11_n_107) & (mul_71_11_n_114 | mul_71_11_n_21));
 assign mul_71_11_n_233 = ~((mul_71_11_n_144 | mul_71_11_n_106) & (mul_71_11_n_123 | mul_71_11_n_21));
 assign mul_71_11_n_232 = ~((mul_71_11_n_144 | mul_71_11_n_116) & (mul_71_11_n_21 | mul_71_11_n_19));
 assign mul_71_11_n_231 = ~((mul_71_11_n_144 | mul_71_11_n_114) & (mul_71_11_n_115 | mul_71_11_n_21));
 assign mul_71_11_n_230 = ~((mul_71_11_n_144 | mul_71_11_n_120) & (mul_71_11_n_118 | mul_71_11_n_21));
 assign mul_71_11_n_229 = ~((mul_71_11_n_144 | mul_71_11_n_110) & (mul_71_11_n_105 | mul_71_11_n_21));
 assign mul_71_11_n_228 = ~((mul_71_11_n_144 | mul_71_11_n_118) & (mul_71_11_n_119 | mul_71_11_n_21));
 assign mul_71_11_n_227 = ~((mul_71_11_n_4 | mul_71_11_n_56) & (mul_71_11_n_81 | mul_71_11_n_55));
 assign mul_71_11_n_226 = ~((mul_71_11_n_4 | mul_71_11_n_42) & (mul_71_11_n_81 | mul_71_11_n_43));
 assign mul_71_11_n_225 = ~((mul_71_11_n_4 | mul_71_11_n_60) & (mul_71_11_n_81 | mul_71_11_n_56));
 assign mul_71_11_n_224 = ~((mul_71_11_n_4 | mul_71_11_n_54) & (mul_71_11_n_81 | mul_71_11_n_61));
 assign mul_71_11_n_223 = ~((mul_71_11_n_4 | mul_71_11_n_46) & (mul_71_11_n_81 | mul_71_11_n_60));
 assign mul_71_11_n_222 = ~((mul_71_11_n_4 | mul_71_11_n_53) & (mul_71_11_n_81 | mul_71_11_n_46));
 assign mul_71_11_n_221 = ~((mul_71_11_n_4 | mul_71_11_n_33) & (mul_71_11_n_81 | mul_71_11_n_48));
 assign mul_71_11_n_220 = ~((mul_71_11_n_4 | mul_71_11_n_45) & (mul_71_11_n_81 | mul_71_11_n_50));
 assign mul_71_11_n_219 = ~((mul_71_11_n_4 | mul_71_11_n_59) & (mul_71_11_n_81 | mul_71_11_n_53));
 assign mul_71_11_n_218 = ~((mul_71_11_n_4 | mul_71_11_n_47) & (mul_71_11_n_81 | mul_71_11_n_52));
 assign mul_71_11_n_217 = ~((mul_71_11_n_4 | mul_71_11_n_50) & (mul_71_11_n_81 | mul_71_11_n_59));
 assign mul_71_11_n_216 = ~((mul_71_11_n_4 | mul_71_11_n_55) & (mul_71_11_n_81 | mul_71_11_n_47));
 assign mul_71_11_n_215 = ~((mul_71_11_n_4 | mul_71_11_n_51) & (mul_71_11_n_81 | mul_71_11_n_58));
 assign mul_71_11_n_214 = ~((mul_71_11_n_4 | mul_71_11_n_52) & (mul_71_11_n_81 | mul_71_11_n_54));
 assign mul_71_11_n_213 = ~((mul_71_11_n_140 | mul_71_11_n_35) & (mul_71_11_n_84 | mul_71_11_n_72));
 assign mul_71_11_n_212 = ~((mul_71_11_n_140 | mul_71_11_n_70) & (mul_71_11_n_84 | mul_71_11_n_127));
 assign mul_71_11_n_211 = ~((mul_71_11_n_140 | mul_71_11_n_100) & (mul_71_11_n_84 | mul_71_11_n_65));
 assign mul_71_11_n_210 = ~((mul_71_11_n_140 | mul_71_11_n_127) & (mul_71_11_n_84 | mul_71_11_n_100));
 assign mul_71_11_n_209 = ~((mul_71_11_n_4 | mul_71_11_n_61) & (mul_71_11_n_81 | mul_71_11_n_51));
 assign mul_71_11_n_208 = ~((mul_71_11_n_140 | mul_71_11_n_41) & (mul_71_11_n_84 | mul_71_11_n_37));
 assign mul_71_11_n_207 = ~((mul_71_11_n_140 | mul_71_11_n_87) & (mul_71_11_n_84 | mul_71_11_n_41));
 assign mul_71_11_n_206 = ~((mul_71_11_n_140 | mul_71_11_n_91) & (mul_71_11_n_84 | mul_71_11_n_62));
 assign mul_71_11_n_205 = ~((mul_71_11_n_4 | mul_71_11_n_58) & (mul_71_11_n_81 | mul_71_11_n_49));
 assign mul_71_11_n_204 = ~((mul_71_11_n_140 | mul_71_11_n_72) & (mul_71_11_n_84 | mul_71_11_n_124));
 assign mul_71_11_n_203 = ~((mul_71_11_n_4 | mul_71_11_n_57) & (mul_71_11_n_81 | mul_71_11_n_45));
 assign mul_71_11_n_202 = ~((mul_71_11_n_140 | mul_71_11_n_124) & (mul_71_11_n_84 | mul_71_11_n_87));
 assign mul_71_11_n_201 = ~((mul_71_11_n_140 | mul_71_11_n_75) & (mul_71_11_n_84 | mul_71_11_n_91));
 assign mul_71_11_n_200 = ((mul_71_11_n_136 & mul_71_11_n_99) | (mul_71_11_n_139 & mul_71_11_n_93));
 assign mul_71_11_n_199 = ~((mul_71_11_n_140 | mul_71_11_n_96) & (mul_71_11_n_84 | mul_71_11_n_75));
 assign mul_71_11_n_198 = ~((mul_71_11_n_140 | mul_71_11_n_65) & (mul_71_11_n_84 | mul_71_11_n_69));
 assign mul_71_11_n_197 = ~((mul_71_11_n_4 | mul_71_11_n_48) & (mul_71_11_n_81 | mul_71_11_n_57));
 assign mul_71_11_n_196 = ~((mul_71_11_n_140 | mul_71_11_n_37) & (mul_71_11_n_84 | mul_71_11_n_38));
 assign mul_71_11_n_195 = ~((mul_71_11_n_140 | mul_71_11_n_97) & (mul_71_11_n_84 | mul_71_11_n_70));
 assign mul_71_11_n_194 = ~((mul_71_11_n_140 | mul_71_11_n_98) & (mul_71_11_n_84 | mul_71_11_n_96));
 assign mul_71_11_n_193 = ~((mul_71_11_n_140 | mul_71_11_n_62) & (mul_71_11_n_84 | mul_71_11_n_92));
 assign mul_71_11_n_192 = ~((mul_71_11_n_140 | mul_71_11_n_38) & (mul_71_11_n_84 | mul_71_11_n_97));
 assign mul_71_11_n_191 = ~((mul_71_11_n_140 | mul_71_11_n_69) & (mul_71_11_n_84 | mul_71_11_n_98));
 assign mul_71_11_n_190 = ~((mul_71_11_n_4 | mul_71_11_n_49) & (mul_71_11_n_81 | mul_71_11_n_42));
 assign mul_71_11_n_189 = ~mul_71_11_n_188;
 assign mul_71_11_n_187 = ~mul_71_11_n_186;
 assign mul_71_11_n_184 = ~((mul_71_11_n_135 | mul_71_11_n_17) & (mul_71_11_n_86 | mul_71_11_n_26));
 assign mul_71_11_n_183 = ~((mul_71_11_n_135 | mul_71_11_n_13) & (mul_71_11_n_86 | mul_71_11_n_27));
 assign mul_71_11_n_182 = ~((mul_71_11_n_135 | mul_71_11_n_10) & (mul_71_11_n_86 | mul_71_11_n_18));
 assign mul_71_11_n_181 = ~((mul_71_11_n_135 | mul_71_11_n_28) & (mul_71_11_n_86 | mul_71_11_n_17));
 assign mul_71_11_n_180 = ~((mul_71_11_n_135 | mul_71_11_n_9) & (mul_71_11_n_86 | mul_71_11_n_11));
 assign mul_71_11_n_179 = ~((mul_71_11_n_135 | mul_71_11_n_14) & (mul_71_11_n_86 | mul_71_11_n_16));
 assign mul_71_11_n_178 = ~((mul_71_11_n_135 | mul_71_11_n_23) & (mul_71_11_n_86 | mul_71_11_n_30));
 assign mul_71_11_n_177 = ~((mul_71_11_n_135 | mul_71_11_n_25) & (mul_71_11_n_86 | mul_71_11_n_14));
 assign mul_71_11_n_176 = ~((mul_71_11_n_135 | mul_71_11_n_29) & (mul_71_11_n_86 | mul_71_11_n_28));
 assign mul_71_11_n_175 = ~((mul_71_11_n_135 | mul_71_11_n_24) & (mul_71_11_n_86 | mul_71_11_n_15));
 assign mul_71_11_n_174 = ~((mul_71_11_n_135 | mul_71_11_n_26) & (mul_71_11_n_86 | mul_71_11_n_24));
 assign mul_71_11_n_173 = ~((mul_71_11_n_135 | mul_71_11_n_8) & (mul_71_11_n_86 | mul_71_11_n_29));
 assign mul_71_11_n_172 = ~((mul_71_11_n_135 | mul_71_11_n_12) & (mul_71_11_n_86 | mul_71_11_n_25));
 assign mul_71_11_n_171 = ~((mul_71_11_n_135 | mul_71_11_n_30) & (mul_71_11_n_86 | mul_71_11_n_12));
 assign mul_71_11_n_170 = ~((mul_71_11_n_135 | mul_71_11_n_18) & (mul_71_11_n_86 | mul_71_11_n_8));
 assign mul_71_11_n_169 = ~((mul_71_11_n_135 | mul_71_11_n_16) & (mul_71_11_n_86 | mul_71_11_n_10));
 assign mul_71_11_n_168 = ~((mul_71_11_n_131 | mul_71_11_n_36) & (mul_71_11_n_83 | mul_71_11_n_94));
 assign mul_71_11_n_167 = ~((mul_71_11_n_131 | mul_71_11_n_77) & (mul_71_11_n_83 | mul_71_11_n_76));
 assign mul_71_11_n_166 = ~((mul_71_11_n_131 | mul_71_11_n_68) & (mul_71_11_n_83 | mul_71_11_n_126));
 assign mul_71_11_n_165 = ~((mul_71_11_n_131 | mul_71_11_n_73) & (mul_71_11_n_83 | mul_71_11_n_88));
 assign mul_71_11_n_164 = ~((mul_71_11_n_131 | mul_71_11_n_71) & (mul_71_11_n_83 | mul_71_11_n_77));
 assign mul_71_11_n_163 = ((mul_71_11_n_82 & mul_71_11_n_74) | (mul_71_11_n_130 & mul_71_11_n_90));
 assign mul_71_11_n_162 = ~((mul_71_11_n_131 | mul_71_11_n_101) & (mul_71_11_n_83 | mul_71_11_n_63));
 assign mul_71_11_n_161 = ~((mul_71_11_n_131 | mul_71_11_n_125) & (mul_71_11_n_83 | mul_71_11_n_71));
 assign mul_71_11_n_160 = ~((mul_71_11_n_131 | mul_71_11_n_67) & (mul_71_11_n_83 | mul_71_11_n_101));
 assign mul_71_11_n_159 = ~((mul_71_11_n_131 | mul_71_11_n_63) & (mul_71_11_n_83 | mul_71_11_n_73));
 assign mul_71_11_n_158 = ~((mul_71_11_n_131 | mul_71_11_n_94) & (mul_71_11_n_83 | mul_71_11_n_95));
 assign mul_71_11_n_157 = ~((mul_71_11_n_131 | mul_71_11_n_66) & (mul_71_11_n_83 | mul_71_11_n_125));
 assign mul_71_11_n_156 = ~((mul_71_11_n_131 | mul_71_11_n_64) & (mul_71_11_n_83 | mul_71_11_n_89));
 assign mul_71_11_n_155 = ~((mul_71_11_n_131 | mul_71_11_n_95) & (mul_71_11_n_83 | mul_71_11_n_67));
 assign mul_71_11_n_154 = ~((mul_71_11_n_131 | mul_71_11_n_39) & (mul_71_11_n_83 | mul_71_11_n_40));
 assign mul_71_11_n_153 = ~((mul_71_11_n_131 | mul_71_11_n_76) & (mul_71_11_n_83 | mul_71_11_n_64));
 assign mul_71_11_n_152 = ~((mul_71_11_n_131 | mul_71_11_n_40) & (mul_71_11_n_83 | mul_71_11_n_68));
 assign mul_71_11_n_151 = ~((mul_71_11_n_131 | mul_71_11_n_126) & (mul_71_11_n_83 | mul_71_11_n_66));
 assign mul_71_11_n_150 = ~((mul_71_11_n_131 | mul_71_11_n_88) & (mul_71_11_n_83 | mul_71_11_n_39));
 assign mul_71_11_n_149 = ~((mul_71_11_n_135 | mul_71_11_n_22) & (mul_71_11_n_86 | mul_71_11_n_23));
 assign mul_71_11_n_148 = ~(mul_71_11_n_134 & n_164);
 assign mul_71_11_n_147 = ~(mul_71_11_n_81 | mul_71_11_n_22);
 assign mul_71_11_n_146 = ~(mul_71_11_n_84 | mul_71_11_n_22);
 assign mul_71_11_n_144 = ~mul_71_11_n_145;
 assign mul_71_11_n_143 = ~mul_71_11_n_4;
 assign mul_71_11_n_142 = ~mul_71_11_n_141;
 assign mul_71_11_n_141 = ~(mul_71_11_n_81 | mul_71_11_n_20);
 assign mul_71_11_n_139 = ~mul_71_11_n_140;
 assign mul_71_11_n_140 = (mul_71_11_n_136 | mul_71_11_n_80);
 assign mul_71_11_n_138 = ~(mul_71_11_n_84 | mul_71_11_n_7);
 assign mul_71_11_n_136 = ~mul_71_11_n_84;
 assign mul_71_11_n_134 = ~mul_71_11_n_135;
 assign mul_71_11_n_133 = ~(mul_71_11_n_86 | mul_71_11_n_22);
 assign mul_71_11_n_132 = ~(mul_71_11_n_83 | mul_71_11_n_22);
 assign mul_71_11_n_130 = ~mul_71_11_n_131;
 assign mul_71_11_n_131 = (mul_71_11_n_82 | mul_71_11_n_79);
 assign mul_71_11_n_129 = ~(mul_71_11_n_83 | mul_71_11_n_6);
 assign mul_71_11_n_122 = ~mul_71_11_n_121;
 assign mul_71_11_n_113 = ~mul_71_11_n_112;
 assign mul_71_11_n_103 = ~mul_71_11_n_102;
 assign mul_71_11_n_93 = ~mul_71_11_n_92;
 assign mul_71_11_n_90 = ~mul_71_11_n_89;
 assign mul_71_11_n_85 = ~mul_71_11_n_86;
 assign mul_71_11_n_82 = ~mul_71_11_n_83;
 assign mul_71_11_n_128 = ({out1[0]} | mul_71_11_n_19);
 assign mul_71_11_n_44 = ~mul_71_11_n_43;
 assign {out1[0]} = ~(mul_71_11_n_21 | mul_71_11_n_22);
 assign mul_71_11_n_27 = ~n_164;
 assign mul_71_11_n_13 = ~n_165;
 assign mul_71_11_n_4 = ~(mul_71_11_n_81 & ~mul_71_11_n_78);
 assign mul_71_11_n_3 = (mul_71_11_n_129 | (mul_71_11_n_130 & mul_71_11_n_74));
endmodule
